-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 4 2021 00:32:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    reset_n_in : in std_logic;
    led_out : out std_logic;
    mosi_in : in std_logic;
    miso_out : out std_logic;
    cs_n_in : in std_logic;
    clk_spi_in : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \GNDG0\ : std_logic;
signal \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net\ : std_logic;
signal \sb_translator_1.cnt_i_0\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \sb_translator_1.cnt_i_1\ : std_logic;
signal \sb_translator_1.cnt19_cry_0\ : std_logic;
signal \sb_translator_1.cnt_RNIOI3OZ0Z_2\ : std_logic;
signal \sb_translator_1.cnt19_cry_1\ : std_logic;
signal \sb_translator_1.cnt_RNISN4OZ0Z_3\ : std_logic;
signal \sb_translator_1.cnt19_cry_2\ : std_logic;
signal \sb_translator_1.cnt_RNI0T5OZ0Z_4\ : std_logic;
signal \sb_translator_1.cnt19_cry_3\ : std_logic;
signal \sb_translator_1.cnt_RNI427OZ0Z_5\ : std_logic;
signal \sb_translator_1.cnt19_cry_4\ : std_logic;
signal \sb_translator_1.cnt_RNI878OZ0Z_6\ : std_logic;
signal \sb_translator_1.cnt19_cry_5\ : std_logic;
signal \sb_translator_1.cnt_RNICC9OZ0Z_7\ : std_logic;
signal \sb_translator_1.cnt19_cry_6\ : std_logic;
signal \sb_translator_1.cnt19_cry_7\ : std_logic;
signal \sb_translator_1.cnt_RNIGHAOZ0Z_8\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \sb_translator_1.cnt_RNIKMBOZ0Z_9\ : std_logic;
signal \sb_translator_1.cnt19_cry_8\ : std_logic;
signal \sb_translator_1.cnt_RNI6O3VZ0Z_10\ : std_logic;
signal \sb_translator_1.cnt19_cry_9\ : std_logic;
signal \sb_translator_1.cnt_RNIO5UPZ0Z_11\ : std_logic;
signal \sb_translator_1.cnt19_cry_10\ : std_logic;
signal \sb_translator_1.cnt_RNISAVPZ0Z_12\ : std_logic;
signal \sb_translator_1.cnt19_cry_11\ : std_logic;
signal \sb_translator_1.cnt_RNI0G0QZ0Z_13\ : std_logic;
signal \sb_translator_1.cnt19_cry_12\ : std_logic;
signal \sb_translator_1.cnt_RNI4L1QZ0Z_14\ : std_logic;
signal \sb_translator_1.cnt19_cry_13\ : std_logic;
signal \sb_translator_1.cnt_RNI8Q2QZ0Z_15\ : std_logic;
signal \sb_translator_1.cnt19_cry_14\ : std_logic;
signal \sb_translator_1.cnt19_cry_15\ : std_logic;
signal \sb_translator_1.cnt_i_16\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \sb_translator_1.cnt19_cry_16\ : std_logic;
signal \sb_translator_1.cnt19_cry_18\ : std_logic;
signal \sb_translator_1.cnt19_cry_20\ : std_logic;
signal \sb_translator_1.cnt19_cry_21\ : std_logic;
signal \sb_translator_1.cnt19_cry_22\ : std_logic;
signal \sb_translator_1.cnt19_cry_23\ : std_logic;
signal \sb_translator_1.cnt19_cry_24\ : std_logic;
signal \sb_translator_1.cnt19_cry_25\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \sb_translator_1.cnt19_cry_26\ : std_logic;
signal \sb_translator_1.cnt19_cry_27\ : std_logic;
signal \sb_translator_1.cnt19_cry_28\ : std_logic;
signal \sb_translator_1.cnt19_cry_29\ : std_logic;
signal \sb_translator_1.cnt19_cry_30\ : std_logic;
signal \sb_translator_1.cnt19_cry_31\ : std_logic;
signal \sb_translator_1.cnt19_cry_32\ : std_logic;
signal \sb_translator_1.cnt19_cry_33\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \sb_translator_1.cnt19_cry_34\ : std_logic;
signal \sb_translator_1.cnt19_cry_35\ : std_logic;
signal \spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4\ : std_logic;
signal \spi_slave_1.un3_mosi_data_out_3\ : std_logic;
signal \spi_slave_1.un3_mosi_data_out_3_cascade_\ : std_logic;
signal \spi_slave_1.bitcnt_rxZ0Z_0\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \spi_slave_1.bitcnt_rxZ0Z_1\ : std_logic;
signal \spi_slave_1.bitcnt_rx_cry_0\ : std_logic;
signal \spi_slave_1.bitcnt_rxZ0Z_2\ : std_logic;
signal \spi_slave_1.bitcnt_rx_cry_1\ : std_logic;
signal \spi_slave_1.bitcnt_rxZ0Z_3\ : std_logic;
signal \spi_slave_1.bitcnt_rx_cry_2\ : std_logic;
signal \spi_slave_1.bitcnt_rx_cry_3\ : std_logic;
signal \spi_slave_1.bitcnt_rxZ0Z_4\ : std_logic;
signal miso_en : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_0\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_1\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_2\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_3\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO\ : std_logic;
signal \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_23\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_18\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_19\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_20\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_21\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_22\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_10\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_2\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_3\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_4\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_5\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_6\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_7\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_8\ : std_logic;
signal \sb_translator_1.stateZ0Z_5\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_13\ : std_logic;
signal \sb_translator_1.cntZ0Z_13\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_14\ : std_logic;
signal \sb_translator_1.cntZ0Z_14\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_15\ : std_logic;
signal \sb_translator_1.cntZ0Z_15\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_16\ : std_logic;
signal \sb_translator_1.cntZ0Z_16\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_1\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_11\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_12\ : std_logic;
signal \sb_translator_1.cnt_RNO_0Z0Z_9\ : std_logic;
signal \sb_translator_1.cntZ0Z_9\ : std_logic;
signal \sb_translator_1.cntZ0Z_12\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_18\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_19\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_20\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_21\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_22\ : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_23\ : std_logic;
signal miso_data_in_19 : std_logic;
signal miso_data_in_20 : std_logic;
signal miso_data_in_21 : std_logic;
signal miso_data_in_22 : std_logic;
signal miso_data_in_23 : std_logic;
signal miso_data_in_8 : std_logic;
signal \spi_slave_1.clk_pos_i\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_22\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_21\ : std_logic;
signal \spi_slave_1.m81_ns_1_cascade_\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_5\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_4\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_20\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_19\ : std_logic;
signal \spi_slave_1.m60_ns_1_cascade_\ : std_logic;
signal clk_spi : std_logic;
signal \spi_slave_1.bitcnt_tx10\ : std_logic;
signal \spi_slave_1.bitcnt_tx10_cascade_\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_8\ : std_logic;
signal miso_tx : std_logic;
signal \spi_slave_1.N_82\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_17\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_10\ : std_logic;
signal \spi_slave_1.m48_ns_1_cascade_\ : std_logic;
signal \spi_slave_1.N_49_0_cascade_\ : std_logic;
signal \spi_slave_1.N_25_0_cascade_\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_23\ : std_logic;
signal \spi_slave_1.miso_data_out_0_sqmuxa\ : std_logic;
signal \spi_slave_1.N_96_mux\ : std_logic;
signal \spi_slave_1.N_94_mux\ : std_logic;
signal \spi_slave_1.N_94_mux_cascade_\ : std_logic;
signal \spi_slave_1.bitcnt_txZ0Z_3\ : std_logic;
signal \spi_slave_1.N_17_0\ : std_logic;
signal \spi_slave_1.N_20_0\ : std_logic;
signal \spi_slave_1.N_91\ : std_logic;
signal miso : std_logic;
signal \spi_slave_1.bitcnt_rxe_0_i\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_1\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_2\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_1\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_3\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_2\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_4\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_3\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_5\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_4\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_6\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_5\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_7\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_6\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_8\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_7\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_8\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_9\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_10\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_9\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_11\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_10\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_12\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_11\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_13\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_12\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_14\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_13\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_15\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_14\ : std_logic;
signal \sb_translator_1.un1_num_leds_0_cry_15\ : std_logic;
signal \sb_translator_1.un1_num_leds_n_16\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_1\ : std_logic;
signal reset_n : std_logic;
signal reset_n_i : std_logic;
signal ram_we_3 : std_logic;
signal ram_we_13 : std_logic;
signal \sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_\ : std_logic;
signal ram_we_5 : std_logic;
signal ram_we_7 : std_logic;
signal ram_we_9 : std_logic;
signal \sb_translator_1.N_1092\ : std_logic;
signal \sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_\ : std_logic;
signal ram_we_11 : std_logic;
signal \sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_\ : std_logic;
signal mosi_data_out_17 : std_logic;
signal demux_data_in_86 : std_logic;
signal demux_data_in_54 : std_logic;
signal \demux.N_877_cascade_\ : std_logic;
signal demux_data_in_70 : std_logic;
signal demux_data_in_62 : std_logic;
signal \demux.N_418_i_0_o2Z0Z_6\ : std_logic;
signal demux_data_in_83 : std_logic;
signal demux_data_in_51 : std_logic;
signal \demux.N_835_cascade_\ : std_logic;
signal demux_data_in_59 : std_logic;
signal demux_data_in_67 : std_logic;
signal \demux.N_421_i_0_o2Z0Z_6\ : std_logic;
signal demux_data_in_63 : std_logic;
signal demux_data_in_57 : std_logic;
signal demux_data_in_87 : std_logic;
signal demux_data_in_79 : std_logic;
signal demux_data_in_55 : std_logic;
signal \demux.N_417_i_0_o2Z0Z_6_cascade_\ : std_logic;
signal \demux.N_890\ : std_logic;
signal demux_data_in_61 : std_logic;
signal demux_data_in_77 : std_logic;
signal demux_data_in_85 : std_logic;
signal demux_data_in_53 : std_logic;
signal \demux.N_419_i_0_o2Z0Z_6_cascade_\ : std_logic;
signal \demux.N_419_i_0_a3Z0Z_1\ : std_logic;
signal demux_data_in_60 : std_logic;
signal demux_data_in_84 : std_logic;
signal demux_data_in_76 : std_logic;
signal demux_data_in_52 : std_logic;
signal \demux.N_420_i_0_o2Z0Z_6_cascade_\ : std_logic;
signal \demux.N_420_i_0_a3Z0Z_1\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_6\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_1\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_3\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_7\ : std_logic;
signal miso_data_in_18 : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_2\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_18\ : std_logic;
signal \spi_slave_1.m72_ns_1\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_14\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_13\ : std_logic;
signal \spi_slave_1.bitcnt_txZ0Z_2\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_12_cascade_\ : std_logic;
signal \spi_slave_1.bitcnt_txZ0Z_1\ : std_logic;
signal \spi_slave_1.m27_ns_1_cascade_\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_7\ : std_logic;
signal \spi_slave_1.N_28_0\ : std_logic;
signal \spi_slave_1.mosi_bufferZ0Z_1\ : std_logic;
signal cs_n : std_logic;
signal mosi : std_logic;
signal \spi_slave_1.mosi_bufferZ0Z_0\ : std_logic;
signal \spi_slave_1.clkZ0Z_0\ : std_logic;
signal \spi_slave_1.clkZ0Z_1\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_17\ : std_logic;
signal \spi_slave_1.bitcnt_rxe_0_i_g\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_9\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_8\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_10\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_11\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_12\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_13\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_14\ : std_logic;
signal mosi_data_out_8 : std_logic;
signal \sb_translator_1.cntZ0Z_0\ : std_logic;
signal mosi_data_out_9 : std_logic;
signal \sb_translator_1.cntZ0Z_1\ : std_logic;
signal \sb_translator_1.cntZ0Z_2\ : std_logic;
signal mosi_data_out_10 : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_16\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_3\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_2\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_5\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_6\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_7\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_4\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_0\ : std_logic;
signal ram_data_in_0 : std_logic;
signal ram_data_in_1 : std_logic;
signal ram_data_in_2 : std_logic;
signal ram_data_in_3 : std_logic;
signal ram_data_in_4 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_5\ : std_logic;
signal mosi_data_out_5 : std_logic;
signal ram_data_in_5 : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_6\ : std_logic;
signal mosi_data_out_6 : std_logic;
signal ram_data_in_6 : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_7\ : std_logic;
signal mosi_data_out_7 : std_logic;
signal ram_data_in_7 : std_logic;
signal ram_we_0 : std_logic;
signal ram_we_2 : std_logic;
signal \sb_translator_1.cnt_RNILAHE_1Z0Z_10\ : std_logic;
signal ram_we_10 : std_logic;
signal ram_we_8 : std_logic;
signal \sb_translator_1.N_1088\ : std_logic;
signal ram_we_12 : std_logic;
signal \sb_translator_1.cnt_RNILAHE_0Z0Z_10\ : std_logic;
signal ram_we_4 : std_logic;
signal \sb_translator_1.cnt_RNIJ7EF_2Z0Z_9\ : std_logic;
signal \sb_translator_1.state_RNI9ILJ_0Z0Z_0\ : std_logic;
signal ram_we_6 : std_logic;
signal \sb_translator_1.cnt_RNIJ7EF_1Z0Z_9\ : std_logic;
signal \sb_translator_1.state_RNI9ILJZ0Z_0\ : std_logic;
signal ram_we_1 : std_logic;
signal \sb_translator_1.N_1091_cascade_\ : std_logic;
signal \sb_translator_1.N_1089_cascade_\ : std_logic;
signal \sb_translator_1.N_1091\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_\ : std_logic;
signal demux_data_in_74 : std_logic;
signal demux_data_in_82 : std_logic;
signal demux_data_in_50 : std_logic;
signal \demux.N_422_i_0_o2Z0Z_6_cascade_\ : std_logic;
signal demux_data_in_73 : std_logic;
signal demux_data_in_81 : std_logic;
signal demux_data_in_49 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_6_cascade_\ : std_logic;
signal \demux.N_423_i_0_a3Z0Z_1\ : std_logic;
signal demux_data_in_58 : std_logic;
signal \demux.N_422_i_0_a3Z0Z_1\ : std_logic;
signal demux_data_in_80 : std_logic;
signal demux_data_in_72 : std_logic;
signal demux_data_in_48 : std_logic;
signal \demux.N_424_i_0_o2_6_cascade_\ : std_logic;
signal demux_data_in_56 : std_logic;
signal \demux.N_424_i_0_a3Z0Z_1\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9\ : std_logic;
signal \sb_translator_1.state_RNIHS98Z0Z_0\ : std_logic;
signal \sb_translator_1.state_RNIHS98_0Z0Z_0\ : std_logic;
signal \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9\ : std_logic;
signal \sb_translator_1.N_1089\ : std_logic;
signal \demux.N_236_cascade_\ : std_logic;
signal \demux.N_235_cascade_\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_6\ : std_logic;
signal ram_sel_6 : std_logic;
signal ram_sel_9 : std_logic;
signal miso_data_in_9 : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_17\ : std_logic;
signal \spi_slave_1.bitcnt_tx_0_sqmuxa\ : std_logic;
signal miso_data_in_10 : std_logic;
signal miso_data_in_11 : std_logic;
signal miso_data_in_12 : std_logic;
signal miso_data_in_13 : std_logic;
signal miso_data_in_14 : std_logic;
signal miso_data_in_15 : std_logic;
signal miso_data_in_16 : std_logic;
signal \sb_translator_1.instr_tmpZ0Z_17\ : std_logic;
signal miso_data_in_17 : std_logic;
signal mosi_data_out_11 : std_logic;
signal \sb_translator_1.cntZ0Z_3\ : std_logic;
signal mosi_data_out_13 : std_logic;
signal \sb_translator_1.cntZ0Z_5\ : std_logic;
signal \sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_9\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_11\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_10\ : std_logic;
signal \sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_\ : std_logic;
signal \sb_translator_1.ram_sel_6_0_0_a2_0_0_7\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10\ : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_0\ : std_logic;
signal addr_out_0 : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_1\ : std_logic;
signal addr_out_1 : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_2\ : std_logic;
signal addr_out_2 : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_3\ : std_logic;
signal addr_out_3 : std_logic;
signal addr_out_4 : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_5\ : std_logic;
signal addr_out_5 : std_logic;
signal addr_out_6 : std_logic;
signal addr_out_7 : std_logic;
signal \sb_translator_1.cnt_RNILAHE_2Z0Z_10\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10\ : std_logic;
signal mosi_data_out_0 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_0\ : std_logic;
signal mosi_data_out_1 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_1\ : std_logic;
signal mosi_data_out_2 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_2\ : std_logic;
signal mosi_data_out_3 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_3\ : std_logic;
signal mosi_data_out_4 : std_logic;
signal \sb_translator_1.instr_tmpZ1Z_4\ : std_logic;
signal \sb_translator_1.state_RNIKJOCZ0Z_5\ : std_logic;
signal \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\ : std_logic;
signal \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11\ : std_logic;
signal \sb_translator_1.cnt19_cry_18_THRU_CO\ : std_logic;
signal \sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_\ : std_logic;
signal mosi_rx : std_logic;
signal \sb_translator_1.state_RNIOH7V9Z0Z_0\ : std_logic;
signal \sb_translator_1.N_58\ : std_logic;
signal \sb_translator_1.state_RNIEL0N9_0Z0Z_6\ : std_logic;
signal \sb_translator_1.cnt_ram_readZ0Z_0\ : std_logic;
signal \sb_translator_1.cnt_ram_readZ0Z_1\ : std_logic;
signal demux_data_in_42 : std_logic;
signal \sb_translator_1.cntZ0Z_11\ : std_logic;
signal \sb_translator_1.cntZ0Z_10\ : std_logic;
signal \sb_translator_1.ram_we_6_0_0_a2_0_6\ : std_logic;
signal miso_data_in_2 : std_logic;
signal mosi_data_out_22 : std_logic;
signal \sb_translator_1.N_1087\ : std_logic;
signal \sb_translator_1.num_leds_1_sqmuxa_cascade_\ : std_logic;
signal \sb_translator_1.send_leds_n_1_sqmuxa\ : std_logic;
signal \sb_translator_1.N_59\ : std_logic;
signal miso_data_in_0 : std_logic;
signal \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5\ : std_logic;
signal \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\ : std_logic;
signal \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0\ : std_logic;
signal mosi_data_out_18 : std_logic;
signal mosi_data_out_19 : std_logic;
signal mosi_data_out_20 : std_logic;
signal \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3\ : std_logic;
signal \demux.N_238_cascade_\ : std_logic;
signal \demux.N_242_cascade_\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_34_cascade_\ : std_logic;
signal \demux.N_424_i_0_aZ0Z2\ : std_logic;
signal \demux.N_242\ : std_logic;
signal \demux.N_916\ : std_logic;
signal ram_sel_5 : std_logic;
signal \demux.N_916_cascade_\ : std_logic;
signal ram_sel_1 : std_logic;
signal \demux.N_239\ : std_logic;
signal \demux.N_241\ : std_logic;
signal \demux.N_915\ : std_logic;
signal ram_sel_12 : std_logic;
signal \demux.N_915_cascade_\ : std_logic;
signal ram_sel_2 : std_logic;
signal ram_sel_3 : std_logic;
signal ram_sel_8 : std_logic;
signal addr_out_8 : std_logic;
signal \sb_translator_1.state_RNI88IGAZ0Z_0\ : std_logic;
signal \sb_translator_1.state_leds_2_sqmuxa\ : std_logic;
signal \sb_translator_1.state_ledsZ0\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_9\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_10\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_13\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_12\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_11\ : std_logic;
signal \spi_slave_1.miso_RNOZ0Z_6\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_16\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_0\ : std_logic;
signal \spi_slave_1.bitcnt_txZ0Z_4\ : std_logic;
signal \spi_slave_1.bitcnt_txZ0Z_0\ : std_logic;
signal \spi_slave_1.N_58_0_cascade_\ : std_logic;
signal \spi_slave_1.miso_data_outZ0Z_15\ : std_logic;
signal \spi_slave_1.N_55_0\ : std_logic;
signal \spi_slave_1.mosi_data_inZ0Z_15\ : std_logic;
signal \spi_slave_1.un3_mosi_data_out_g\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_5\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_6\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_7\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_8\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_3\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_4\ : std_logic;
signal \sb_translator_1.cnt19\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_2\ : std_logic;
signal \sb_translator_1.state56_a_5_44_cascade_\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_1\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_0\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_1\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_0\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_2\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_1\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_3\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_2\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_4\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_3\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_5\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_4\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_6\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_5\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_7\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_6\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_7\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_8\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_8\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_10\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_9\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_11\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_10\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_11\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_12\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_13\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_14\ : std_logic;
signal \sb_translator_1.cnt_leds_cry_15\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1\ : std_logic;
signal demux_data_in_40 : std_logic;
signal demux_data_in_88 : std_logic;
signal \demux.N_424_i_0_a3Z0Z_4\ : std_logic;
signal demux_data_in_8 : std_logic;
signal \demux.N_424_i_0_o2Z0Z_1_cascade_\ : std_logic;
signal demux_data_in_0 : std_logic;
signal \demux.N_424_i_0_aZ0Z3_cascade_\ : std_logic;
signal demux_data_in_35 : std_logic;
signal demux_data_in_107 : std_logic;
signal demux_data_in_91 : std_logic;
signal \demux.N_421_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_2 : std_logic;
signal demux_data_in_106 : std_logic;
signal demux_data_in_34 : std_logic;
signal \demux.N_422_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_90 : std_logic;
signal \demux.N_422_i_0_a3Z0Z_4\ : std_logic;
signal demux_data_in_10 : std_logic;
signal \demux.N_422_i_0_o2Z0Z_1_cascade_\ : std_logic;
signal demux_data_in_9 : std_logic;
signal demux_data_in_89 : std_logic;
signal \demux.N_423_i_0_a3Z0Z_5_cascade_\ : std_logic;
signal demux_data_in_43 : std_logic;
signal \demux.N_837\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_34\ : std_logic;
signal \demux.N_918_cascade_\ : std_logic;
signal demux_data_in_105 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_5_cascade_\ : std_logic;
signal demux_data_in_33 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_0\ : std_logic;
signal \demux.N_918\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_7\ : std_logic;
signal \demux.N_424_i_0_o2_0_1\ : std_logic;
signal \demux.N_236\ : std_logic;
signal \demux.N_235\ : std_logic;
signal \demux.N_424_i_0_o2_0Z0Z_2\ : std_logic;
signal \demux.N_237\ : std_logic;
signal \demux.N_424_i_0_o2_0_8Z0Z_1_cascade_\ : std_logic;
signal \demux.N_238\ : std_logic;
signal \demux.N_917\ : std_logic;
signal \demux.N_424_i_0_o2_0_7_cascade_\ : std_logic;
signal \demux.N_424_i_0_o2_0_10\ : std_logic;
signal \demux.N_424_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_16 : std_logic;
signal demux_data_in_96 : std_logic;
signal demux_data_in_64 : std_logic;
signal \demux.N_424_i_0_o2Z0Z_4_cascade_\ : std_logic;
signal \demux.N_424_i_0_o2Z0Z_8\ : std_logic;
signal \demux.N_424_i_0_aZ0Z3\ : std_logic;
signal \demux.N_424_i_0_o2_9\ : std_logic;
signal \demux.N_424_i_0_o2Z0Z_8_cascade_\ : std_logic;
signal \demux.N_424_i_0_o2Z0Z_7\ : std_logic;
signal demux_data_in_24 : std_logic;
signal \demux.N_424_i_0_a3Z0Z_7\ : std_logic;
signal ram_sel_0 : std_logic;
signal ram_sel_11 : std_logic;
signal \demux.N_906_cascade_\ : std_logic;
signal ram_sel_4 : std_logic;
signal \demux.N_424_i_0_o2_0Z0Z_3\ : std_logic;
signal demux_data_in_28 : std_logic;
signal ram_sel_13 : std_logic;
signal ram_sel_10 : std_logic;
signal ram_sel_7 : std_logic;
signal \demux.N_240\ : std_logic;
signal demux_data_in_29 : std_logic;
signal \sb_translator_1.state56_a_5_ac0_1\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIJDTTZ0Z_2\ : std_logic;
signal \sb_translator_1.state56_a_5_44\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_0_c_THRU_CO\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIPJTTZ0Z_3\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_0\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIERUEZ0Z_3\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIVPTTZ0Z_4\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_1\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIHUUEZ0Z_4\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI50UTZ0Z_5\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_2\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIB6UTZ0Z_6\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_3\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIHCUTZ0Z_7\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_4\ : std_logic;
signal \sb_translator_1.cnt_leds_RNINIUTZ0Z_8\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_5\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_6\ : std_logic;
signal \sb_translator_1.num_leds_RNITOUTZ0Z_8\ : std_logic;
signal \sb_translator_1.cnt_leds_RNITAVEZ0Z_8\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \sb_translator_1.num_leds_RNIH2E91Z0Z_9\ : std_logic;
signal \sb_translator_1.num_leds_RNI0EVEZ0Z_8\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_7\ : std_logic;
signal \sb_translator_1.num_leds_RNICJVN1Z0Z_10\ : std_logic;
signal \sb_translator_1.num_leds_RNIHKEQZ0Z_9\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_8\ : std_logic;
signal \sb_translator_1.num_leds_RNIP02R1Z0Z_11\ : std_logic;
signal \sb_translator_1.num_leds_RNIRUGTZ0Z_10\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_9\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_10\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_11\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_12\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_13\ : std_logic;
signal \sb_translator_1.state56_a_5_cry_14\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_16\ : std_logic;
signal \sb_translator_1.cnt_leds_i_16_cascade_\ : std_logic;
signal \sb_translator_1.num_leds_RNIOJBMZ0Z_15\ : std_logic;
signal \sb_translator_1.num_leds_RNIU1HTZ0Z_11\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIV62R1Z0Z_13\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI48HTZ0Z_14\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_15\ : std_logic;
signal \sb_translator_1.cnt_leds_i_16\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_15\ : std_logic;
signal \sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_12\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_13\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI15HTZ0Z_13\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_14\ : std_logic;
signal \sb_translator_1.num_ledsZ0Z_13\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_14\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14\ : std_logic;
signal demux_data_in_66 : std_logic;
signal demux_data_in_30 : std_logic;
signal demux_data_in_102 : std_logic;
signal demux_data_in_32 : std_logic;
signal demux_data_in_104 : std_logic;
signal \demux.N_424_i_0_o2_0Z0Z_0\ : std_logic;
signal demux_data_in_44 : std_logic;
signal demux_data_in_22 : std_logic;
signal \demux.N_418_i_0_o2Z0Z_4\ : std_logic;
signal demux_data_in_78 : std_logic;
signal \demux.N_884_cascade_\ : std_logic;
signal demux_data_in_27 : std_logic;
signal demux_data_in_19 : std_logic;
signal demux_data_in_99 : std_logic;
signal demux_data_in_75 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_0\ : std_logic;
signal \demux.N_421_i_0_o2Z0Z_4_cascade_\ : std_logic;
signal \demux.N_421_i_0_a3Z0Z_7\ : std_logic;
signal demux_data_in_11 : std_logic;
signal \demux.N_421_i_0_o2Z0Z_8_cascade_\ : std_logic;
signal \demux.N_421_i_0_o2Z0Z_2\ : std_logic;
signal \demux.N_422_i_0_o2Z0Z_8\ : std_logic;
signal \demux.N_422_i_0_o2Z0Z_9\ : std_logic;
signal \demux.N_422_i_0_aZ0Z3\ : std_logic;
signal \demux.N_422_i_0_o2Z0Z_7\ : std_logic;
signal \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1\ : std_logic;
signal mosi_data_out_16 : std_logic;
signal \sb_translator_1.cntZ0Z_8\ : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_8\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_12\ : std_logic;
signal \sb_translator_1.cnt_ledsZ0Z_9\ : std_logic;
signal \sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9\ : std_logic;
signal demux_data_in_26 : std_logic;
signal \demux.N_422_i_0_a3Z0Z_7\ : std_logic;
signal demux_data_in_15 : std_logic;
signal demux_data_in_25 : std_logic;
signal demux_data_in_17 : std_logic;
signal demux_data_in_97 : std_logic;
signal demux_data_in_65 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_4_cascade_\ : std_logic;
signal \demux.N_423_i_0_a3Z0Z_7\ : std_logic;
signal demux_data_in_41 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_8_cascade_\ : std_logic;
signal \demux.N_423_i_0_o2Z0Z_2\ : std_logic;
signal demux_data_in_111 : std_logic;
signal demux_data_in_39 : std_logic;
signal demux_data_in_95 : std_logic;
signal \demux.N_417_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal \demux.N_417_i_0_o2Z0Z_1\ : std_logic;
signal demux_data_in_47 : std_logic;
signal \demux.N_417_i_0_a3Z0Z_4\ : std_logic;
signal demux_data_in_109 : std_logic;
signal demux_data_in_37 : std_logic;
signal demux_data_in_93 : std_logic;
signal \demux.N_419_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_45 : std_logic;
signal \demux.N_419_i_0_o2Z0Z_2_cascade_\ : std_logic;
signal demux_data_in_13 : std_logic;
signal \demux.N_419_i_0_a3Z0Z_5\ : std_logic;
signal demux_data_in_69 : std_logic;
signal \demux.N_419_i_0_a3Z0Z_7\ : std_logic;
signal \demux.N_419_i_0_o2Z0Z_8\ : std_logic;
signal \sb_translator_1.state56_a_5_6\ : std_logic;
signal \sb_translator_1.state56_a_5_11\ : std_logic;
signal \sb_translator_1.state56_a_5_5\ : std_logic;
signal \sb_translator_1.state56_a_5_13\ : std_logic;
signal \sb_translator_1.state56_a_5_14\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_12_cascade_\ : std_logic;
signal \sb_translator_1.state56_17\ : std_logic;
signal \sb_translator_1.state_leds_RNIGMAHZ0\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_15_cascade_\ : std_logic;
signal \sb_translator_1.N_712_cascade_\ : std_logic;
signal \sb_translator_1.num_leds_1_sqmuxa\ : std_logic;
signal \sb_translator_1.stateZ0Z_7\ : std_logic;
signal \sb_translator_1.state56_a_5_2\ : std_logic;
signal \sb_translator_1.state56_a_5_7\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_0\ : std_logic;
signal \sb_translator_1.state56_a_5_12\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_8\ : std_logic;
signal \sb_translator_1.N_729\ : std_logic;
signal \sb_translator_1.N_712\ : std_logic;
signal \sb_translator_1.stateZ0Z_0\ : std_logic;
signal \sb_translator_1.state_RNIOCIR9Z0Z_5\ : std_logic;
signal \sb_translator_1.state56_a_5_4\ : std_logic;
signal \sb_translator_1.state56_a_5_10\ : std_logic;
signal \sb_translator_1.state56_a_5_3\ : std_logic;
signal \sb_translator_1.state56_a_5_16\ : std_logic;
signal \sb_translator_1.state56_a_5_8\ : std_logic;
signal \sb_translator_1.state56_a_5_9\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_11_cascade_\ : std_logic;
signal \sb_translator_1.state56_a_5_15\ : std_logic;
signal \sb_translator_1.N_318_i_i_o2_14\ : std_logic;
signal \sb_translator_1.state_RNII30CZ0Z_0\ : std_logic;
signal \sb_translator_1.stateZ0Z_1\ : std_logic;
signal mosi_data_out_23 : std_logic;
signal mosi_data_out_21 : std_logic;
signal \sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0\ : std_logic;
signal mosi_data_out_12 : std_logic;
signal \sb_translator_1.cntZ0Z_4\ : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_4\ : std_logic;
signal mosi_data_out_14 : std_logic;
signal \sb_translator_1.cntZ0Z_6\ : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_6\ : std_logic;
signal \sb_translator_1.stateZ0Z_6\ : std_logic;
signal mosi_data_out_15 : std_logic;
signal \sb_translator_1.cntZ0Z_7\ : std_logic;
signal \sb_translator_1.addr_out_RNO_0Z0Z_7\ : std_logic;
signal \ws2812.new_data_req_e_1\ : std_logic;
signal \ws2812.N_140_cascade_\ : std_logic;
signal ws2812_next_led : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_0\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_10\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_12\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_18\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_15\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_16\ : std_logic;
signal demux_data_in_94 : std_logic;
signal demux_data_in_110 : std_logic;
signal \demux.N_418_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_38 : std_logic;
signal demux_data_in_46 : std_logic;
signal \demux.N_418_i_0_o2Z0Z_1_cascade_\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_8\ : std_logic;
signal demux_data_in_14 : std_logic;
signal \demux.N_880\ : std_logic;
signal demux_data_in_36 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_4\ : std_logic;
signal \demux.N_424_i_0_a2Z0Z_5\ : std_logic;
signal demux_data_in_108 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_11\ : std_logic;
signal \demux.N_420_i_0_o2Z0Z_0_cascade_\ : std_logic;
signal demux_data_in_92 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_2\ : std_logic;
signal demux_data_in_12 : std_logic;
signal \demux.N_420_i_0_o2Z0Z_1_cascade_\ : std_logic;
signal \demux.N_420_i_0_a3Z0Z_4\ : std_logic;
signal demux_data_in_7 : std_logic;
signal \demux.N_888_cascade_\ : std_logic;
signal demux_data_in_6 : std_logic;
signal \demux.N_874_cascade_\ : std_logic;
signal demux_data_in_4 : std_logic;
signal \demux.N_417_i_0_o2Z0Z_9\ : std_logic;
signal \demux.N_888\ : std_logic;
signal \demux.N_417_i_0_o2Z0Z_7\ : std_logic;
signal miso_data_in_7 : std_logic;
signal \demux.N_874\ : std_logic;
signal \demux.N_418_i_0_o2Z0Z_8\ : std_logic;
signal \demux.N_418_i_0_o2Z0Z_9\ : std_logic;
signal \demux.N_418_i_0_o2Z0Z_7\ : std_logic;
signal miso_data_in_6 : std_logic;
signal miso_data_in_5 : std_logic;
signal \demux.N_421_i_0_o2Z0Z_9\ : std_logic;
signal demux_data_in_3 : std_logic;
signal \demux.N_421_i_0_o2Z0Z_10\ : std_logic;
signal miso_data_in_3 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_9\ : std_logic;
signal demux_data_in_1 : std_logic;
signal \demux.N_423_i_0_o2Z0Z_10\ : std_logic;
signal miso_data_in_1 : std_logic;
signal miso_data_in_4 : std_logic;
signal \sb_translator_1.state_g_1\ : std_logic;
signal demux_data_in_31 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_1\ : std_logic;
signal demux_data_in_71 : std_logic;
signal \demux.N_417_i_0_a3Z0Z_7_cascade_\ : std_logic;
signal \demux.N_417_i_0_o2Z0Z_8\ : std_logic;
signal demux_data_in_103 : std_logic;
signal demux_data_in_23 : std_logic;
signal \demux.N_417_i_0_o2Z0Z_4\ : std_logic;
signal demux_data_in_18 : std_logic;
signal demux_data_in_98 : std_logic;
signal \demux.N_422_i_0_o2Z0Z_4\ : std_logic;
signal demux_data_in_101 : std_logic;
signal demux_data_in_21 : std_logic;
signal \demux.N_419_i_0_o2Z0Z_4\ : std_logic;
signal demux_data_in_100 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_3\ : std_logic;
signal demux_data_in_20 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_10\ : std_logic;
signal demux_data_in_68 : std_logic;
signal \demux.N_424_i_0_a2Z0Z_9\ : std_logic;
signal \demux.N_420_i_0_o2Z0Z_4_cascade_\ : std_logic;
signal \demux.N_420_i_0_a3Z0Z_7\ : std_logic;
signal \ws2812.state_ns_0_i_o2_6_0_cascade_\ : std_logic;
signal \ws2812.N_105_cascade_\ : std_logic;
signal \ws2812.state_ns_0_i_o2_6_0\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \ws2812.bit_counter_RNI5NQB3Z0Z_1\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_0\ : std_logic;
signal \ws2812.bit_counter_0_RNIJC643Z0Z_0\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_1\ : std_logic;
signal \ws2812.bit_counterZ0Z_3\ : std_logic;
signal \ws2812.bit_counter_0_RNIKD643Z0Z_1\ : std_logic;
signal \ws2812.bit_counter_0_RNO_0Z0Z_1\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_2\ : std_logic;
signal \ws2812.bit_counter_0_RNILE643Z0Z_2\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_3\ : std_logic;
signal \ws2812.bit_counter_0_RNIMF643Z0Z_3\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_4\ : std_logic;
signal \ws2812.bit_counter_RNI6OQB3Z0Z_2\ : std_logic;
signal \ws2812.bit_counter_6\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_5\ : std_logic;
signal \ws2812.bit_counter_RNI7PQB3Z0Z_3\ : std_logic;
signal \ws2812.bit_counter_7\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_6\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_7\ : std_logic;
signal \ws2812.bit_counter_RNI8QQB3Z0Z_4\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \ws2812.bit_counter_RNI9RQB3Z0Z_5\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_8\ : std_logic;
signal \ws2812.bit_counter_0_RNING643Z0Z_4\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_9\ : std_logic;
signal \ws2812.un1_bit_counter_12_axb_11\ : std_logic;
signal \ws2812.un1_bit_counter_12_cry_10\ : std_logic;
signal \ws2812.state_ns_0_i_o2_7_0\ : std_logic;
signal \ws2812.bit_counterZ0Z_4\ : std_logic;
signal \ws2812.bit_counterZ0Z_5\ : std_logic;
signal \ws2812.bit_counter_8\ : std_logic;
signal \ws2812.N_52_cascade_\ : std_logic;
signal led : std_logic;
signal rgb_data_out_12 : std_logic;
signal rgb_data_out_15 : std_logic;
signal rgb_data_out_10 : std_logic;
signal \ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_\ : std_logic;
signal \ws2812.rgb_counter_RNI2H7OZ0Z_2\ : std_logic;
signal \ws2812.rgb_counter_RNIFI3MZ0Z_2\ : std_logic;
signal \ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_\ : std_logic;
signal \ws2812.N_108_cascade_\ : std_logic;
signal \ws2812.N_107\ : std_logic;
signal \ws2812.rgb_counter_RNI4J7OZ0Z_2\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_8\ : std_logic;
signal rgb_data_out_8 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_13\ : std_logic;
signal rgb_data_out_13 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_11\ : std_logic;
signal rgb_data_out_11 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_9\ : std_logic;
signal rgb_data_out_9 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_1\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_21\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_20\ : std_logic;
signal \sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1\ : std_logic;
signal \demux.N_424_i_0_o2Z0Z_0\ : std_logic;
signal \demux.N_419_i_0_o2Z0Z_9\ : std_logic;
signal demux_data_in_5 : std_logic;
signal \demux.N_419_i_0_o2Z0Z_10\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_5\ : std_logic;
signal \demux.N_420_i_0_o2Z0Z_8\ : std_logic;
signal \demux.N_420_i_0_o2Z0Z_9\ : std_logic;
signal \demux.N_420_i_0_aZ0Z3\ : std_logic;
signal \demux.N_420_i_0_o2Z0Z_7\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_4\ : std_logic;
signal \sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1\ : std_logic;
signal \ws2812.stateZ0Z_1\ : std_logic;
signal \ws2812.state_ns_0_i_o2_8_0\ : std_logic;
signal \ws2812.bit_counterZ0Z_1\ : std_logic;
signal \ws2812.bit_counterZ0Z_0\ : std_logic;
signal \ws2812.bit_counter_11\ : std_logic;
signal \ws2812.bit_counter_0_RNO_0Z0Z_4\ : std_logic;
signal \ws2812.bit_counter_0_RNO_0Z0Z_0\ : std_logic;
signal \ws2812.bit_counterZ0Z_2\ : std_logic;
signal \ws2812.bit_counter_i_0\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \ws2812.un6_data_axb_1\ : std_logic;
signal \ws2812.un6_data_cry_0\ : std_logic;
signal \ws2812.bit_counter_0_RNIQAT2Z0Z_0\ : std_logic;
signal \ws2812.un6_data_cry_1\ : std_logic;
signal \ws2812.bit_counter_0_RNIRBT2Z0Z_1\ : std_logic;
signal \ws2812.un6_data_cry_2\ : std_logic;
signal \ws2812.bit_counter_0_RNISCT2Z0Z_2\ : std_logic;
signal \ws2812.un6_data_cry_3_c_RNIKNFBZ0\ : std_logic;
signal \ws2812.un6_data_cry_3\ : std_logic;
signal \ws2812.bit_counter_0_RNITDT2Z0Z_3\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ws2812.un6_data_cry_4_c_RNIMQGBZ0\ : std_logic;
signal \ws2812.un6_data_cry_4\ : std_logic;
signal \ws2812.un6_data_axb_6\ : std_logic;
signal \ws2812.un6_data_cry_5\ : std_logic;
signal \ws2812.un6_data_axb_7\ : std_logic;
signal \ws2812.un6_data_cry_6\ : std_logic;
signal \ws2812.un6_data_cry_7\ : std_logic;
signal \ws2812.un6_data_axb_8\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \ws2812.un6_data_cry_8\ : std_logic;
signal \ws2812.un6_data_cry_9\ : std_logic;
signal \ws2812.un6_data_axb_11\ : std_logic;
signal \ws2812.un6_data_cry_10\ : std_logic;
signal \ws2812.data_RNOZ0Z_11\ : std_logic;
signal \ws2812.data_RNOZ0Z_12\ : std_logic;
signal \ws2812.data_RNOZ0Z_13\ : std_logic;
signal \ws2812.un6_data_cry_11\ : std_logic;
signal \ws2812.bit_counter_10\ : std_logic;
signal \ws2812.un6_data_axb_10\ : std_logic;
signal \ws2812.bit_counter_9\ : std_logic;
signal \ws2812.un6_data_axb_9\ : std_logic;
signal \ws2812.data_RNOZ0Z_6\ : std_logic;
signal \ws2812.data_RNOZ0Z_5\ : std_logic;
signal \ws2812.data_5_iv_0_47_a2_0_a2_0\ : std_logic;
signal \ws2812.data_5_iv_0_47_a2_0_a2_6_1\ : std_logic;
signal \ws2812.data_5_iv_0_47_a2_0_a2_6\ : std_logic;
signal \ws2812.data_RNOZ0Z_10\ : std_logic;
signal \ws2812.data_RNOZ0Z_9\ : std_logic;
signal \ws2812.data_RNOZ0Z_8\ : std_logic;
signal \ws2812.N_135\ : std_logic;
signal \ws2812.data_RNOZ0Z_2\ : std_logic;
signal \ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_\ : std_logic;
signal \ws2812.N_115\ : std_logic;
signal rgb_data_out_16 : std_logic;
signal rgb_data_out_0 : std_logic;
signal rgb_data_out_20 : std_logic;
signal \ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_\ : std_logic;
signal rgb_data_out_4 : std_logic;
signal \ws2812.N_127\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \ws2812.un1_rgb_counter_cry_0\ : std_logic;
signal \ws2812.un1_rgb_counter_cry_1\ : std_logic;
signal \ws2812.rgb_counter_RNO_0Z0Z_3\ : std_logic;
signal \ws2812.un1_rgb_counter_cry_2\ : std_logic;
signal \ws2812.un1_rgb_counter_cry_3\ : std_logic;
signal rgb_data_out_1 : std_logic;
signal rgb_data_out_21 : std_logic;
signal \ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_\ : std_logic;
signal rgb_data_out_5 : std_logic;
signal \ws2812.N_120\ : std_logic;
signal rgb_data_out_18 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_2\ : std_logic;
signal rgb_data_out_2 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_17\ : std_logic;
signal rgb_data_out_17 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_23\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_14\ : std_logic;
signal rgb_data_out_14 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_22\ : std_logic;
signal \ws2812.N_105\ : std_logic;
signal rgb_data_out_23 : std_logic;
signal \ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_\ : std_logic;
signal \ws2812.N_117\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_3\ : std_logic;
signal rgb_data_out_3 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_19\ : std_logic;
signal rgb_data_out_19 : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_7\ : std_logic;
signal rgb_data_out_7 : std_logic;
signal \ws2812.rgb_counter_4\ : std_logic;
signal rgb_data_out_22 : std_logic;
signal \ws2812.rgb_data_pmux_6_i_m2_ns_1\ : std_logic;
signal \ws2812.N_124\ : std_logic;
signal \ws2812.rgb_counter_0_sqmuxa_0_a2_0_1\ : std_logic;
signal \ws2812.rgb_counterZ0Z_2\ : std_logic;
signal \ws2812.rgb_counter_RNI2AOD3Z0Z_2\ : std_logic;
signal \ws2812.rgb_counterZ0Z_1\ : std_logic;
signal \ws2812.rgb_counter_RNI19OD3Z0Z_1\ : std_logic;
signal \ws2812.rgb_counterZ0Z_3\ : std_logic;
signal \ws2812.rgb_counter_RNI3BOD3Z0Z_3\ : std_logic;
signal \ws2812.rgb_counterZ0Z_0\ : std_logic;
signal \ws2812.un1_rgb_counter_cry_0_c_RNOZ0\ : std_logic;
signal \ws2812.N_106\ : std_logic;
signal send_leds_n : std_logic;
signal \ws2812.stateZ0Z_0\ : std_logic;
signal \ws2812.N_228\ : std_logic;
signal \ws2812.state_RNIELS35Z0Z_0\ : std_logic;
signal \sb_translator_1.rgb_data_tmpZ0Z_6\ : std_logic;
signal rgb_data_out_6 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_sb : std_logic;
signal \sb_translator_1.state_leds_2_sqmuxa_g\ : std_logic;
signal reset_n_i_g : std_logic;

signal reset_n_in_wire : std_logic;
signal clk_spi_in_wire : std_logic;
signal miso_out_wire : std_logic;
signal cs_n_in_wire : std_logic;
signal mosi_in_wire : std_logic;
signal led_out_wire : std_logic;
signal \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    reset_n_in_wire <= reset_n_in;
    clk_spi_in_wire <= clk_spi_in;
    miso_out <= miso_out_wire;
    cs_n_in_wire <= cs_n_in;
    mosi_in_wire <= mosi_in;
    led_out <= led_out_wire;
    demux_data_in_15 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_14 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_13 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_12 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_11 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_10 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_9 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_8 <= \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18112\&\N__16216\&\N__16432\&\N__16633\&\N__14785\&\N__15004\&\N__15232\&\N__15451\&\N__15655\;
    \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18115\&\N__16210\&\N__16426\&\N__16660\&\N__14788\&\N__15013\&\N__15259\&\N__15454\&\N__15688\;
    \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13492\&'0'&\N__13671\&'0'&\N__13818\&'0'&\N__12641\&'0'&\N__12753\&'0'&\N__12909\&'0'&\N__13028\&'0'&\N__13143\;
    demux_data_in_23 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_22 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_21 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_20 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_19 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_18 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_17 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_16 <= \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18088\&\N__16192\&\N__16408\&\N__16609\&\N__14760\&\N__14980\&\N__15208\&\N__15427\&\N__15631\;
    \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18091\&\N__16186\&\N__16402\&\N__16636\&\N__14763\&\N__14989\&\N__15235\&\N__15430\&\N__15664\;
    \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13471\&'0'&\N__13672\&'0'&\N__13830\&'0'&\N__12653\&'0'&\N__12776\&'0'&\N__12910\&'0'&\N__13029\&'0'&\N__13144\;
    demux_data_in_87 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_86 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_85 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_84 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_83 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_82 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_81 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_80 <= \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18208\&\N__16310\&\N__16526\&\N__16727\&\N__14881\&\N__15100\&\N__15326\&\N__15547\&\N__15751\;
    \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18211\&\N__16306\&\N__16522\&\N__16744\&\N__14884\&\N__15109\&\N__15343\&\N__15550\&\N__15777\;
    \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13491\&'0'&\N__13670\&'0'&\N__13798\&'0'&\N__12654\&'0'&\N__12757\&'0'&\N__12906\&'0'&\N__13024\&'0'&\N__13152\;
    demux_data_in_47 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_46 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_45 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_44 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_43 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_42 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_41 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_40 <= \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18178\&\N__16261\&\N__16477\&\N__16678\&\N__14863\&\N__15091\&\N__15277\&\N__15505\&\N__15718\;
    \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18181\&\N__16279\&\N__16495\&\N__16699\&\N__14878\&\N__15082\&\N__15298\&\N__15508\&\N__15745\;
    \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13440\&'0'&\N__13611\&'0'&\N__13788\&'0'&\N__12635\&'0'&\N__12692\&'0'&\N__12856\&'0'&\N__12948\&'0'&\N__13070\;
    demux_data_in_95 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_94 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_93 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_92 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_91 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_90 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_89 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_88 <= \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18184\&\N__16288\&\N__16504\&\N__16705\&\N__14857\&\N__15076\&\N__15304\&\N__15523\&\N__15727\;
    \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18187\&\N__16282\&\N__16498\&\N__16730\&\N__14860\&\N__15085\&\N__15329\&\N__15526\&\N__15760\;
    \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13472\&'0'&\N__13645\&'0'&\N__13789\&'0'&\N__12642\&'0'&\N__12775\&'0'&\N__12907\&'0'&\N__12977\&'0'&\N__13098\;
    demux_data_in_7 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_6 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_5 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_4 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_3 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_2 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_1 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_0 <= \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18228\&\N__16324\&\N__16540\&\N__16743\&\N__14905\&\N__15124\&\N__15342\&\N__15561\&\N__15773\;
    \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18229\&\N__16323\&\N__16539\&\N__16750\&\N__14906\&\N__15129\&\N__15349\&\N__15562\&\N__15784\;
    \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13487\&'0'&\N__13669\&'0'&\N__13822\&'0'&\N__12655\&'0'&\N__12777\&'0'&\N__12896\&'0'&\N__13030\&'0'&\N__13156\;
    demux_data_in_39 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_38 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_37 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_36 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_35 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_34 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_33 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_32 <= \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18202\&\N__16285\&\N__16501\&\N__16702\&\N__14887\&\N__15115\&\N__15301\&\N__15529\&\N__15742\;
    \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18205\&\N__16303\&\N__16519\&\N__16723\&\N__14902\&\N__15106\&\N__15322\&\N__15532\&\N__15767\;
    \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13460\&'0'&\N__13634\&'0'&\N__13823\&'0'&\N__12636\&'0'&\N__12771\&'0'&\N__12873\&'0'&\N__12986\&'0'&\N__13107\;
    demux_data_in_55 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_54 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_53 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_52 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_51 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_50 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_49 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_48 <= \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18154\&\N__16237\&\N__16453\&\N__16654\&\N__14839\&\N__15067\&\N__15253\&\N__15481\&\N__15694\;
    \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18157\&\N__16255\&\N__16471\&\N__16675\&\N__14854\&\N__15058\&\N__15274\&\N__15484\&\N__15721\;
    \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13450\&'0'&\N__13624\&'0'&\N__13802\&'0'&\N__12630\&'0'&\N__12761\&'0'&\N__12866\&'0'&\N__12978\&'0'&\N__13099\;
    demux_data_in_31 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_30 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_29 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_28 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_27 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_26 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_25 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_24 <= \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18226\&\N__16309\&\N__16525\&\N__16726\&\N__14907\&\N__15130\&\N__15325\&\N__15553\&\N__15766\;
    \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18227\&\N__16322\&\N__16538\&\N__16742\&\N__14911\&\N__15128\&\N__15341\&\N__15554\&\N__15780\;
    \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13484\&'0'&\N__13662\&'0'&\N__13824\&'0'&\N__12652\&'0'&\N__12783\&'0'&\N__12897\&'0'&\N__13009\&'0'&\N__13127\;
    demux_data_in_111 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_110 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_109 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_108 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_107 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_106 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_105 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_104 <= \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18136\&\N__16240\&\N__16456\&\N__16657\&\N__14809\&\N__15028\&\N__15256\&\N__15475\&\N__15679\;
    \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18139\&\N__16234\&\N__16450\&\N__16684\&\N__14812\&\N__15037\&\N__15283\&\N__15478\&\N__15712\;
    \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13476\&'0'&\N__13665\&'0'&\N__13791\&'0'&\N__12640\&'0'&\N__12752\&'0'&\N__12905\&'0'&\N__13011\&'0'&\N__13145\;
    demux_data_in_103 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_102 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_101 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_100 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_99 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_98 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_97 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_96 <= \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18160\&\N__16264\&\N__16480\&\N__16681\&\N__14833\&\N__15052\&\N__15280\&\N__15499\&\N__15703\;
    \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18163\&\N__16258\&\N__16474\&\N__16708\&\N__14836\&\N__15061\&\N__15307\&\N__15502\&\N__15736\;
    \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13477\&'0'&\N__13655\&'0'&\N__13790\&'0'&\N__12643\&'0'&\N__12751\&'0'&\N__12904\&'0'&\N__13010\&'0'&\N__13128\;
    demux_data_in_63 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_62 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_61 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_60 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_59 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_58 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_57 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_56 <= \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18130\&\N__16213\&\N__16429\&\N__16630\&\N__14815\&\N__15043\&\N__15229\&\N__15457\&\N__15670\;
    \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18133\&\N__16231\&\N__16447\&\N__16651\&\N__14830\&\N__15034\&\N__15250\&\N__15460\&\N__15697\;
    \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13464\&'0'&\N__13638\&'0'&\N__13825\&'0'&\N__12631\&'0'&\N__12778\&'0'&\N__12895\&'0'&\N__12979\&'0'&\N__13100\;
    demux_data_in_71 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_70 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_69 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_68 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_67 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_66 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_65 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_64 <= \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18106\&\N__16189\&\N__16405\&\N__16606\&\N__14791\&\N__15019\&\N__15205\&\N__15433\&\N__15646\;
    \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18109\&\N__16207\&\N__16423\&\N__16627\&\N__14806\&\N__15010\&\N__15226\&\N__15436\&\N__15673\;
    \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13485\&'0'&\N__13663\&'0'&\N__13826\&'0'&\N__12650\&'0'&\N__12779\&'0'&\N__12894\&'0'&\N__13007\&'0'&\N__13125\;
    demux_data_in_79 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(14);
    demux_data_in_78 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(12);
    demux_data_in_77 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(10);
    demux_data_in_76 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(8);
    demux_data_in_75 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(6);
    demux_data_in_74 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(4);
    demux_data_in_73 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(2);
    demux_data_in_72 <= \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\(0);
    \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__18082\&\N__16164\&\N__16380\&\N__16581\&\N__14766\&\N__14995\&\N__15180\&\N__15409\&\N__15622\;
    \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__18085\&\N__16183\&\N__16399\&\N__16603\&\N__14782\&\N__14986\&\N__15202\&\N__15412\&\N__15649\;
    \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__13486\&'0'&\N__13664\&'0'&\N__13831\&'0'&\N__12651\&'0'&\N__12784\&'0'&\N__12908\&'0'&\N__13008\&'0'&\N__13126\;

    \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26207\,
            WCLKE => \N__13897\,
            WCLK => \N__27513\,
            WE => \N__26214\
        );

    \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26212\,
            WCLKE => \N__13324\,
            WCLK => \N__27520\,
            WE => \N__26218\
        );

    \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26156\,
            WCLKE => \N__13288\,
            WCLK => \N__27463\,
            WE => \N__26170\
        );

    \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26066\,
            WCLKE => \N__11197\,
            WCLK => \N__27431\,
            WE => \N__26125\
        );

    \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26172\,
            WCLKE => \N__11353\,
            WCLK => \N__27478\,
            WE => \N__26196\
        );

    \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26155\,
            WCLKE => \N__13339\,
            WCLK => \N__27447\,
            WE => \N__26097\
        );

    \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__25951\,
            WCLKE => \N__14035\,
            WCLK => \N__27424\,
            WE => \N__26034\
        );

    \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26177\,
            WCLKE => \N__13969\,
            WCLK => \N__27443\,
            WE => \N__26078\
        );

    \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__25949\,
            WCLKE => \N__11230\,
            WCLK => \N__27420\,
            WE => \N__25950\
        );

    \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26191\,
            WCLKE => \N__11215\,
            WCLK => \N__27503\,
            WE => \N__26213\
        );

    \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26173\,
            WCLKE => \N__13237\,
            WCLK => \N__27492\,
            WE => \N__26197\
        );

    \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26178\,
            WCLKE => \N__11191\,
            WCLK => \N__27455\,
            WE => \N__26148\
        );

    \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26153\,
            WCLKE => \N__13270\,
            WCLK => \N__27473\,
            WE => \N__26149\
        );

    \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net\,
            RE => \N__26154\,
            WCLKE => \N__11173\,
            WCLK => \N__27488\,
            WE => \N__26195\
        );

    \reset_n_input_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__28196\,
            DIN => \N__28195\,
            DOUT => \N__28194\,
            PACKAGEPIN => reset_n_in_wire
        );

    \reset_n_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28196\,
            PADOUT => \N__28195\,
            PADIN => \N__28194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => reset_n,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_spi_input_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__28187\,
            DIN => \N__28186\,
            DOUT => \N__28185\,
            PACKAGEPIN => clk_spi_in_wire
        );

    \clk_spi_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28187\,
            PADOUT => \N__28186\,
            PADIN => \N__28185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_spi,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \miso_output_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__28178\,
            DIN => \N__28177\,
            DOUT => \N__28176\,
            PACKAGEPIN => miso_out_wire
        );

    \miso_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28178\,
            PADOUT => \N__28177\,
            PADIN => \N__28176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \cs_n_input_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__28169\,
            DIN => \N__28168\,
            DOUT => \N__28167\,
            PACKAGEPIN => cs_n_in_wire
        );

    \cs_n_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28169\,
            PADOUT => \N__28168\,
            PADIN => \N__28167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => cs_n,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \mosi_input_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__28160\,
            DIN => \N__28159\,
            DOUT => \N__28158\,
            PACKAGEPIN => mosi_in_wire
        );

    \mosi_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28160\,
            PADOUT => \N__28159\,
            PADIN => \N__28158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => mosi,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__28151\,
            DIN => \N__28150\,
            DOUT => \N__28149\,
            PACKAGEPIN => led_out_wire
        );

    \led_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__28151\,
            PADOUT => \N__28150\,
            PADIN => \N__28149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24811\,
            INPUTCLK => \GNDG0\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6847\ : CascadeMux
    port map (
            O => \N__28132\,
            I => \N__28129\
        );

    \I__6846\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28126\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__28126\,
            I => \ws2812.rgb_counter_0_sqmuxa_0_a2_0_1\
        );

    \I__6844\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28119\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__28122\,
            I => \N__28103\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28100\
        );

    \I__6841\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28097\
        );

    \I__6840\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28088\
        );

    \I__6839\ : InMux
    port map (
            O => \N__28116\,
            I => \N__28088\
        );

    \I__6838\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28088\
        );

    \I__6837\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28088\
        );

    \I__6836\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28083\
        );

    \I__6835\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28083\
        );

    \I__6834\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28078\
        );

    \I__6833\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28078\
        );

    \I__6832\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28073\
        );

    \I__6831\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28073\
        );

    \I__6830\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28068\
        );

    \I__6829\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28068\
        );

    \I__6828\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28065\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__28100\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__28097\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__28088\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__28083\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__28078\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__28073\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__28068\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__28065\,
            I => \ws2812.rgb_counterZ0Z_2\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__6818\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28042\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__28042\,
            I => \ws2812.rgb_counter_RNI2AOD3Z0Z_2\
        );

    \I__6816\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28036\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28029\
        );

    \I__6814\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28026\
        );

    \I__6813\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28023\
        );

    \I__6812\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28020\
        );

    \I__6811\ : InMux
    port map (
            O => \N__28032\,
            I => \N__28017\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__28029\,
            I => \ws2812.rgb_counterZ0Z_1\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__28026\,
            I => \ws2812.rgb_counterZ0Z_1\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__28023\,
            I => \ws2812.rgb_counterZ0Z_1\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__28020\,
            I => \ws2812.rgb_counterZ0Z_1\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__28017\,
            I => \ws2812.rgb_counterZ0Z_1\
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__28006\,
            I => \N__28003\
        );

    \I__6804\ : InMux
    port map (
            O => \N__28003\,
            I => \N__28000\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__28000\,
            I => \ws2812.rgb_counter_RNI19OD3Z0Z_1\
        );

    \I__6802\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27991\
        );

    \I__6801\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27988\
        );

    \I__6800\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27985\
        );

    \I__6799\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27982\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__27991\,
            I => \N__27979\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27976\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27973\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27970\
        );

    \I__6794\ : Span4Mux_v
    port map (
            O => \N__27979\,
            I => \N__27967\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__27976\,
            I => \N__27964\
        );

    \I__6792\ : Span4Mux_s3_h
    port map (
            O => \N__27973\,
            I => \N__27961\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__27970\,
            I => \N__27958\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__27967\,
            I => \ws2812.rgb_counterZ0Z_3\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__27964\,
            I => \ws2812.rgb_counterZ0Z_3\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__27961\,
            I => \ws2812.rgb_counterZ0Z_3\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__27958\,
            I => \ws2812.rgb_counterZ0Z_3\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__27949\,
            I => \N__27946\
        );

    \I__6785\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27943\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__27943\,
            I => \ws2812.rgb_counter_RNI3BOD3Z0Z_3\
        );

    \I__6783\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27928\
        );

    \I__6781\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27925\
        );

    \I__6780\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27922\
        );

    \I__6779\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27917\
        );

    \I__6778\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27917\
        );

    \I__6777\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27912\
        );

    \I__6776\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27912\
        );

    \I__6775\ : Span4Mux_v
    port map (
            O => \N__27928\,
            I => \N__27908\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__27925\,
            I => \N__27903\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__27922\,
            I => \N__27903\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__27917\,
            I => \N__27900\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__27912\,
            I => \N__27897\
        );

    \I__6770\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27894\
        );

    \I__6769\ : Span4Mux_s0_h
    port map (
            O => \N__27908\,
            I => \N__27889\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__27903\,
            I => \N__27889\
        );

    \I__6767\ : Span4Mux_v
    port map (
            O => \N__27900\,
            I => \N__27886\
        );

    \I__6766\ : Span4Mux_s3_h
    port map (
            O => \N__27897\,
            I => \N__27883\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__27894\,
            I => \ws2812.rgb_counterZ0Z_0\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__27889\,
            I => \ws2812.rgb_counterZ0Z_0\
        );

    \I__6763\ : Odrv4
    port map (
            O => \N__27886\,
            I => \ws2812.rgb_counterZ0Z_0\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__27883\,
            I => \ws2812.rgb_counterZ0Z_0\
        );

    \I__6761\ : CascadeMux
    port map (
            O => \N__27874\,
            I => \N__27871\
        );

    \I__6760\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27868\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__27868\,
            I => \ws2812.un1_rgb_counter_cry_0_c_RNOZ0\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__27865\,
            I => \N__27852\
        );

    \I__6757\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27845\
        );

    \I__6756\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27845\
        );

    \I__6755\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27845\
        );

    \I__6754\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27842\
        );

    \I__6753\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27831\
        );

    \I__6752\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27831\
        );

    \I__6751\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27831\
        );

    \I__6750\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27831\
        );

    \I__6749\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27831\
        );

    \I__6748\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27825\
        );

    \I__6747\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27822\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__27845\,
            I => \N__27819\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__27842\,
            I => \N__27814\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27814\
        );

    \I__6743\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27809\
        );

    \I__6742\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27809\
        );

    \I__6741\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27806\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27801\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27801\
        );

    \I__6738\ : Span4Mux_v
    port map (
            O => \N__27819\,
            I => \N__27796\
        );

    \I__6737\ : Span4Mux_v
    port map (
            O => \N__27814\,
            I => \N__27796\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__27809\,
            I => \ws2812.N_106\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__27806\,
            I => \ws2812.N_106\
        );

    \I__6734\ : Odrv12
    port map (
            O => \N__27801\,
            I => \ws2812.N_106\
        );

    \I__6733\ : Odrv4
    port map (
            O => \N__27796\,
            I => \ws2812.N_106\
        );

    \I__6732\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27783\
        );

    \I__6731\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27780\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27777\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__27780\,
            I => \N__27774\
        );

    \I__6728\ : Span4Mux_s0_h
    port map (
            O => \N__27777\,
            I => \N__27771\
        );

    \I__6727\ : Span12Mux_s7_v
    port map (
            O => \N__27774\,
            I => \N__27766\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__27771\,
            I => \N__27763\
        );

    \I__6725\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27758\
        );

    \I__6724\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27758\
        );

    \I__6723\ : Odrv12
    port map (
            O => \N__27766\,
            I => send_leds_n
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__27763\,
            I => send_leds_n
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__27758\,
            I => send_leds_n
        );

    \I__6720\ : CascadeMux
    port map (
            O => \N__27751\,
            I => \N__27738\
        );

    \I__6719\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27727\
        );

    \I__6718\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27727\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__27748\,
            I => \N__27724\
        );

    \I__6716\ : CascadeMux
    port map (
            O => \N__27747\,
            I => \N__27720\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__27746\,
            I => \N__27716\
        );

    \I__6714\ : CascadeMux
    port map (
            O => \N__27745\,
            I => \N__27712\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__27744\,
            I => \N__27708\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27705\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__27742\,
            I => \N__27702\
        );

    \I__6710\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27697\
        );

    \I__6709\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27693\
        );

    \I__6708\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27680\
        );

    \I__6707\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27680\
        );

    \I__6706\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27680\
        );

    \I__6705\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27680\
        );

    \I__6704\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27680\
        );

    \I__6703\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27680\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__27727\,
            I => \N__27676\
        );

    \I__6701\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27661\
        );

    \I__6700\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27661\
        );

    \I__6699\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27661\
        );

    \I__6698\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27661\
        );

    \I__6697\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27661\
        );

    \I__6696\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27661\
        );

    \I__6695\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27661\
        );

    \I__6694\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27658\
        );

    \I__6693\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27647\
        );

    \I__6692\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27647\
        );

    \I__6691\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27647\
        );

    \I__6690\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27647\
        );

    \I__6689\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27647\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27644\
        );

    \I__6687\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27641\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__27693\,
            I => \N__27636\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27636\
        );

    \I__6684\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27633\
        );

    \I__6683\ : Span12Mux_s5_v
    port map (
            O => \N__27676\,
            I => \N__27628\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__27661\,
            I => \N__27628\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__27658\,
            I => \N__27621\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27621\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__27644\,
            I => \N__27621\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__27641\,
            I => \N__27616\
        );

    \I__6677\ : Span4Mux_h
    port map (
            O => \N__27636\,
            I => \N__27616\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__27633\,
            I => \ws2812.stateZ0Z_0\
        );

    \I__6675\ : Odrv12
    port map (
            O => \N__27628\,
            I => \ws2812.stateZ0Z_0\
        );

    \I__6674\ : Odrv4
    port map (
            O => \N__27621\,
            I => \ws2812.stateZ0Z_0\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__27616\,
            I => \ws2812.stateZ0Z_0\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__27607\,
            I => \N__27604\
        );

    \I__6671\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27601\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27597\
        );

    \I__6669\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27594\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__27597\,
            I => \N__27589\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27589\
        );

    \I__6666\ : Span4Mux_h
    port map (
            O => \N__27589\,
            I => \N__27585\
        );

    \I__6665\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27582\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__27585\,
            I => \ws2812.N_228\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__27582\,
            I => \ws2812.N_228\
        );

    \I__6662\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27569\
        );

    \I__6661\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27569\
        );

    \I__6660\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27566\
        );

    \I__6659\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27563\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27559\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__27566\,
            I => \N__27556\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__27563\,
            I => \N__27553\
        );

    \I__6655\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27550\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__27559\,
            I => \N__27545\
        );

    \I__6653\ : Span4Mux_h
    port map (
            O => \N__27556\,
            I => \N__27545\
        );

    \I__6652\ : Span4Mux_h
    port map (
            O => \N__27553\,
            I => \N__27540\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__27550\,
            I => \N__27540\
        );

    \I__6650\ : Odrv4
    port map (
            O => \N__27545\,
            I => \ws2812.state_RNIELS35Z0Z_0\
        );

    \I__6649\ : Odrv4
    port map (
            O => \N__27540\,
            I => \ws2812.state_RNIELS35Z0Z_0\
        );

    \I__6648\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27532\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27529\
        );

    \I__6646\ : Odrv12
    port map (
            O => \N__27529\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_6\
        );

    \I__6645\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27523\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__27523\,
            I => rgb_data_out_6
        );

    \I__6643\ : ClkMux
    port map (
            O => \N__27520\,
            I => \N__27214\
        );

    \I__6642\ : ClkMux
    port map (
            O => \N__27519\,
            I => \N__27214\
        );

    \I__6641\ : ClkMux
    port map (
            O => \N__27518\,
            I => \N__27214\
        );

    \I__6640\ : ClkMux
    port map (
            O => \N__27517\,
            I => \N__27214\
        );

    \I__6639\ : ClkMux
    port map (
            O => \N__27516\,
            I => \N__27214\
        );

    \I__6638\ : ClkMux
    port map (
            O => \N__27515\,
            I => \N__27214\
        );

    \I__6637\ : ClkMux
    port map (
            O => \N__27514\,
            I => \N__27214\
        );

    \I__6636\ : ClkMux
    port map (
            O => \N__27513\,
            I => \N__27214\
        );

    \I__6635\ : ClkMux
    port map (
            O => \N__27512\,
            I => \N__27214\
        );

    \I__6634\ : ClkMux
    port map (
            O => \N__27511\,
            I => \N__27214\
        );

    \I__6633\ : ClkMux
    port map (
            O => \N__27510\,
            I => \N__27214\
        );

    \I__6632\ : ClkMux
    port map (
            O => \N__27509\,
            I => \N__27214\
        );

    \I__6631\ : ClkMux
    port map (
            O => \N__27508\,
            I => \N__27214\
        );

    \I__6630\ : ClkMux
    port map (
            O => \N__27507\,
            I => \N__27214\
        );

    \I__6629\ : ClkMux
    port map (
            O => \N__27506\,
            I => \N__27214\
        );

    \I__6628\ : ClkMux
    port map (
            O => \N__27505\,
            I => \N__27214\
        );

    \I__6627\ : ClkMux
    port map (
            O => \N__27504\,
            I => \N__27214\
        );

    \I__6626\ : ClkMux
    port map (
            O => \N__27503\,
            I => \N__27214\
        );

    \I__6625\ : ClkMux
    port map (
            O => \N__27502\,
            I => \N__27214\
        );

    \I__6624\ : ClkMux
    port map (
            O => \N__27501\,
            I => \N__27214\
        );

    \I__6623\ : ClkMux
    port map (
            O => \N__27500\,
            I => \N__27214\
        );

    \I__6622\ : ClkMux
    port map (
            O => \N__27499\,
            I => \N__27214\
        );

    \I__6621\ : ClkMux
    port map (
            O => \N__27498\,
            I => \N__27214\
        );

    \I__6620\ : ClkMux
    port map (
            O => \N__27497\,
            I => \N__27214\
        );

    \I__6619\ : ClkMux
    port map (
            O => \N__27496\,
            I => \N__27214\
        );

    \I__6618\ : ClkMux
    port map (
            O => \N__27495\,
            I => \N__27214\
        );

    \I__6617\ : ClkMux
    port map (
            O => \N__27494\,
            I => \N__27214\
        );

    \I__6616\ : ClkMux
    port map (
            O => \N__27493\,
            I => \N__27214\
        );

    \I__6615\ : ClkMux
    port map (
            O => \N__27492\,
            I => \N__27214\
        );

    \I__6614\ : ClkMux
    port map (
            O => \N__27491\,
            I => \N__27214\
        );

    \I__6613\ : ClkMux
    port map (
            O => \N__27490\,
            I => \N__27214\
        );

    \I__6612\ : ClkMux
    port map (
            O => \N__27489\,
            I => \N__27214\
        );

    \I__6611\ : ClkMux
    port map (
            O => \N__27488\,
            I => \N__27214\
        );

    \I__6610\ : ClkMux
    port map (
            O => \N__27487\,
            I => \N__27214\
        );

    \I__6609\ : ClkMux
    port map (
            O => \N__27486\,
            I => \N__27214\
        );

    \I__6608\ : ClkMux
    port map (
            O => \N__27485\,
            I => \N__27214\
        );

    \I__6607\ : ClkMux
    port map (
            O => \N__27484\,
            I => \N__27214\
        );

    \I__6606\ : ClkMux
    port map (
            O => \N__27483\,
            I => \N__27214\
        );

    \I__6605\ : ClkMux
    port map (
            O => \N__27482\,
            I => \N__27214\
        );

    \I__6604\ : ClkMux
    port map (
            O => \N__27481\,
            I => \N__27214\
        );

    \I__6603\ : ClkMux
    port map (
            O => \N__27480\,
            I => \N__27214\
        );

    \I__6602\ : ClkMux
    port map (
            O => \N__27479\,
            I => \N__27214\
        );

    \I__6601\ : ClkMux
    port map (
            O => \N__27478\,
            I => \N__27214\
        );

    \I__6600\ : ClkMux
    port map (
            O => \N__27477\,
            I => \N__27214\
        );

    \I__6599\ : ClkMux
    port map (
            O => \N__27476\,
            I => \N__27214\
        );

    \I__6598\ : ClkMux
    port map (
            O => \N__27475\,
            I => \N__27214\
        );

    \I__6597\ : ClkMux
    port map (
            O => \N__27474\,
            I => \N__27214\
        );

    \I__6596\ : ClkMux
    port map (
            O => \N__27473\,
            I => \N__27214\
        );

    \I__6595\ : ClkMux
    port map (
            O => \N__27472\,
            I => \N__27214\
        );

    \I__6594\ : ClkMux
    port map (
            O => \N__27471\,
            I => \N__27214\
        );

    \I__6593\ : ClkMux
    port map (
            O => \N__27470\,
            I => \N__27214\
        );

    \I__6592\ : ClkMux
    port map (
            O => \N__27469\,
            I => \N__27214\
        );

    \I__6591\ : ClkMux
    port map (
            O => \N__27468\,
            I => \N__27214\
        );

    \I__6590\ : ClkMux
    port map (
            O => \N__27467\,
            I => \N__27214\
        );

    \I__6589\ : ClkMux
    port map (
            O => \N__27466\,
            I => \N__27214\
        );

    \I__6588\ : ClkMux
    port map (
            O => \N__27465\,
            I => \N__27214\
        );

    \I__6587\ : ClkMux
    port map (
            O => \N__27464\,
            I => \N__27214\
        );

    \I__6586\ : ClkMux
    port map (
            O => \N__27463\,
            I => \N__27214\
        );

    \I__6585\ : ClkMux
    port map (
            O => \N__27462\,
            I => \N__27214\
        );

    \I__6584\ : ClkMux
    port map (
            O => \N__27461\,
            I => \N__27214\
        );

    \I__6583\ : ClkMux
    port map (
            O => \N__27460\,
            I => \N__27214\
        );

    \I__6582\ : ClkMux
    port map (
            O => \N__27459\,
            I => \N__27214\
        );

    \I__6581\ : ClkMux
    port map (
            O => \N__27458\,
            I => \N__27214\
        );

    \I__6580\ : ClkMux
    port map (
            O => \N__27457\,
            I => \N__27214\
        );

    \I__6579\ : ClkMux
    port map (
            O => \N__27456\,
            I => \N__27214\
        );

    \I__6578\ : ClkMux
    port map (
            O => \N__27455\,
            I => \N__27214\
        );

    \I__6577\ : ClkMux
    port map (
            O => \N__27454\,
            I => \N__27214\
        );

    \I__6576\ : ClkMux
    port map (
            O => \N__27453\,
            I => \N__27214\
        );

    \I__6575\ : ClkMux
    port map (
            O => \N__27452\,
            I => \N__27214\
        );

    \I__6574\ : ClkMux
    port map (
            O => \N__27451\,
            I => \N__27214\
        );

    \I__6573\ : ClkMux
    port map (
            O => \N__27450\,
            I => \N__27214\
        );

    \I__6572\ : ClkMux
    port map (
            O => \N__27449\,
            I => \N__27214\
        );

    \I__6571\ : ClkMux
    port map (
            O => \N__27448\,
            I => \N__27214\
        );

    \I__6570\ : ClkMux
    port map (
            O => \N__27447\,
            I => \N__27214\
        );

    \I__6569\ : ClkMux
    port map (
            O => \N__27446\,
            I => \N__27214\
        );

    \I__6568\ : ClkMux
    port map (
            O => \N__27445\,
            I => \N__27214\
        );

    \I__6567\ : ClkMux
    port map (
            O => \N__27444\,
            I => \N__27214\
        );

    \I__6566\ : ClkMux
    port map (
            O => \N__27443\,
            I => \N__27214\
        );

    \I__6565\ : ClkMux
    port map (
            O => \N__27442\,
            I => \N__27214\
        );

    \I__6564\ : ClkMux
    port map (
            O => \N__27441\,
            I => \N__27214\
        );

    \I__6563\ : ClkMux
    port map (
            O => \N__27440\,
            I => \N__27214\
        );

    \I__6562\ : ClkMux
    port map (
            O => \N__27439\,
            I => \N__27214\
        );

    \I__6561\ : ClkMux
    port map (
            O => \N__27438\,
            I => \N__27214\
        );

    \I__6560\ : ClkMux
    port map (
            O => \N__27437\,
            I => \N__27214\
        );

    \I__6559\ : ClkMux
    port map (
            O => \N__27436\,
            I => \N__27214\
        );

    \I__6558\ : ClkMux
    port map (
            O => \N__27435\,
            I => \N__27214\
        );

    \I__6557\ : ClkMux
    port map (
            O => \N__27434\,
            I => \N__27214\
        );

    \I__6556\ : ClkMux
    port map (
            O => \N__27433\,
            I => \N__27214\
        );

    \I__6555\ : ClkMux
    port map (
            O => \N__27432\,
            I => \N__27214\
        );

    \I__6554\ : ClkMux
    port map (
            O => \N__27431\,
            I => \N__27214\
        );

    \I__6553\ : ClkMux
    port map (
            O => \N__27430\,
            I => \N__27214\
        );

    \I__6552\ : ClkMux
    port map (
            O => \N__27429\,
            I => \N__27214\
        );

    \I__6551\ : ClkMux
    port map (
            O => \N__27428\,
            I => \N__27214\
        );

    \I__6550\ : ClkMux
    port map (
            O => \N__27427\,
            I => \N__27214\
        );

    \I__6549\ : ClkMux
    port map (
            O => \N__27426\,
            I => \N__27214\
        );

    \I__6548\ : ClkMux
    port map (
            O => \N__27425\,
            I => \N__27214\
        );

    \I__6547\ : ClkMux
    port map (
            O => \N__27424\,
            I => \N__27214\
        );

    \I__6546\ : ClkMux
    port map (
            O => \N__27423\,
            I => \N__27214\
        );

    \I__6545\ : ClkMux
    port map (
            O => \N__27422\,
            I => \N__27214\
        );

    \I__6544\ : ClkMux
    port map (
            O => \N__27421\,
            I => \N__27214\
        );

    \I__6543\ : ClkMux
    port map (
            O => \N__27420\,
            I => \N__27214\
        );

    \I__6542\ : ClkMux
    port map (
            O => \N__27419\,
            I => \N__27214\
        );

    \I__6541\ : GlobalMux
    port map (
            O => \N__27214\,
            I => \N__27211\
        );

    \I__6540\ : DummyBuf
    port map (
            O => \N__27211\,
            I => clk_sb
        );

    \I__6539\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27201\
        );

    \I__6538\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27201\
        );

    \I__6537\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27198\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27188\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__27198\,
            I => \N__27185\
        );

    \I__6534\ : CEMux
    port map (
            O => \N__27197\,
            I => \N__27166\
        );

    \I__6533\ : CEMux
    port map (
            O => \N__27196\,
            I => \N__27166\
        );

    \I__6532\ : CEMux
    port map (
            O => \N__27195\,
            I => \N__27166\
        );

    \I__6531\ : CEMux
    port map (
            O => \N__27194\,
            I => \N__27166\
        );

    \I__6530\ : CEMux
    port map (
            O => \N__27193\,
            I => \N__27166\
        );

    \I__6529\ : CEMux
    port map (
            O => \N__27192\,
            I => \N__27166\
        );

    \I__6528\ : CEMux
    port map (
            O => \N__27191\,
            I => \N__27166\
        );

    \I__6527\ : Glb2LocalMux
    port map (
            O => \N__27188\,
            I => \N__27166\
        );

    \I__6526\ : Glb2LocalMux
    port map (
            O => \N__27185\,
            I => \N__27166\
        );

    \I__6525\ : GlobalMux
    port map (
            O => \N__27166\,
            I => \N__27163\
        );

    \I__6524\ : gio2CtrlBuf
    port map (
            O => \N__27163\,
            I => \sb_translator_1.state_leds_2_sqmuxa_g\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__27160\,
            I => \N__27154\
        );

    \I__6522\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27150\
        );

    \I__6521\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27143\
        );

    \I__6520\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27143\
        );

    \I__6519\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27143\
        );

    \I__6518\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27140\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27120\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__27143\,
            I => \N__27117\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27104\
        );

    \I__6514\ : SRMux
    port map (
            O => \N__27139\,
            I => \N__26920\
        );

    \I__6513\ : SRMux
    port map (
            O => \N__27138\,
            I => \N__26920\
        );

    \I__6512\ : SRMux
    port map (
            O => \N__27137\,
            I => \N__26920\
        );

    \I__6511\ : SRMux
    port map (
            O => \N__27136\,
            I => \N__26920\
        );

    \I__6510\ : SRMux
    port map (
            O => \N__27135\,
            I => \N__26920\
        );

    \I__6509\ : SRMux
    port map (
            O => \N__27134\,
            I => \N__26920\
        );

    \I__6508\ : SRMux
    port map (
            O => \N__27133\,
            I => \N__26920\
        );

    \I__6507\ : SRMux
    port map (
            O => \N__27132\,
            I => \N__26920\
        );

    \I__6506\ : SRMux
    port map (
            O => \N__27131\,
            I => \N__26920\
        );

    \I__6505\ : SRMux
    port map (
            O => \N__27130\,
            I => \N__26920\
        );

    \I__6504\ : SRMux
    port map (
            O => \N__27129\,
            I => \N__26920\
        );

    \I__6503\ : SRMux
    port map (
            O => \N__27128\,
            I => \N__26920\
        );

    \I__6502\ : SRMux
    port map (
            O => \N__27127\,
            I => \N__26920\
        );

    \I__6501\ : SRMux
    port map (
            O => \N__27126\,
            I => \N__26920\
        );

    \I__6500\ : SRMux
    port map (
            O => \N__27125\,
            I => \N__26920\
        );

    \I__6499\ : SRMux
    port map (
            O => \N__27124\,
            I => \N__26920\
        );

    \I__6498\ : SRMux
    port map (
            O => \N__27123\,
            I => \N__26920\
        );

    \I__6497\ : Glb2LocalMux
    port map (
            O => \N__27120\,
            I => \N__26920\
        );

    \I__6496\ : Glb2LocalMux
    port map (
            O => \N__27117\,
            I => \N__26920\
        );

    \I__6495\ : SRMux
    port map (
            O => \N__27116\,
            I => \N__26920\
        );

    \I__6494\ : SRMux
    port map (
            O => \N__27115\,
            I => \N__26920\
        );

    \I__6493\ : SRMux
    port map (
            O => \N__27114\,
            I => \N__26920\
        );

    \I__6492\ : SRMux
    port map (
            O => \N__27113\,
            I => \N__26920\
        );

    \I__6491\ : SRMux
    port map (
            O => \N__27112\,
            I => \N__26920\
        );

    \I__6490\ : SRMux
    port map (
            O => \N__27111\,
            I => \N__26920\
        );

    \I__6489\ : SRMux
    port map (
            O => \N__27110\,
            I => \N__26920\
        );

    \I__6488\ : SRMux
    port map (
            O => \N__27109\,
            I => \N__26920\
        );

    \I__6487\ : SRMux
    port map (
            O => \N__27108\,
            I => \N__26920\
        );

    \I__6486\ : SRMux
    port map (
            O => \N__27107\,
            I => \N__26920\
        );

    \I__6485\ : Glb2LocalMux
    port map (
            O => \N__27104\,
            I => \N__26920\
        );

    \I__6484\ : SRMux
    port map (
            O => \N__27103\,
            I => \N__26920\
        );

    \I__6483\ : SRMux
    port map (
            O => \N__27102\,
            I => \N__26920\
        );

    \I__6482\ : SRMux
    port map (
            O => \N__27101\,
            I => \N__26920\
        );

    \I__6481\ : SRMux
    port map (
            O => \N__27100\,
            I => \N__26920\
        );

    \I__6480\ : SRMux
    port map (
            O => \N__27099\,
            I => \N__26920\
        );

    \I__6479\ : SRMux
    port map (
            O => \N__27098\,
            I => \N__26920\
        );

    \I__6478\ : SRMux
    port map (
            O => \N__27097\,
            I => \N__26920\
        );

    \I__6477\ : SRMux
    port map (
            O => \N__27096\,
            I => \N__26920\
        );

    \I__6476\ : SRMux
    port map (
            O => \N__27095\,
            I => \N__26920\
        );

    \I__6475\ : SRMux
    port map (
            O => \N__27094\,
            I => \N__26920\
        );

    \I__6474\ : SRMux
    port map (
            O => \N__27093\,
            I => \N__26920\
        );

    \I__6473\ : SRMux
    port map (
            O => \N__27092\,
            I => \N__26920\
        );

    \I__6472\ : SRMux
    port map (
            O => \N__27091\,
            I => \N__26920\
        );

    \I__6471\ : SRMux
    port map (
            O => \N__27090\,
            I => \N__26920\
        );

    \I__6470\ : SRMux
    port map (
            O => \N__27089\,
            I => \N__26920\
        );

    \I__6469\ : SRMux
    port map (
            O => \N__27088\,
            I => \N__26920\
        );

    \I__6468\ : SRMux
    port map (
            O => \N__27087\,
            I => \N__26920\
        );

    \I__6467\ : SRMux
    port map (
            O => \N__27086\,
            I => \N__26920\
        );

    \I__6466\ : SRMux
    port map (
            O => \N__27085\,
            I => \N__26920\
        );

    \I__6465\ : SRMux
    port map (
            O => \N__27084\,
            I => \N__26920\
        );

    \I__6464\ : SRMux
    port map (
            O => \N__27083\,
            I => \N__26920\
        );

    \I__6463\ : SRMux
    port map (
            O => \N__27082\,
            I => \N__26920\
        );

    \I__6462\ : SRMux
    port map (
            O => \N__27081\,
            I => \N__26920\
        );

    \I__6461\ : SRMux
    port map (
            O => \N__27080\,
            I => \N__26920\
        );

    \I__6460\ : SRMux
    port map (
            O => \N__27079\,
            I => \N__26920\
        );

    \I__6459\ : SRMux
    port map (
            O => \N__27078\,
            I => \N__26920\
        );

    \I__6458\ : SRMux
    port map (
            O => \N__27077\,
            I => \N__26920\
        );

    \I__6457\ : SRMux
    port map (
            O => \N__27076\,
            I => \N__26920\
        );

    \I__6456\ : SRMux
    port map (
            O => \N__27075\,
            I => \N__26920\
        );

    \I__6455\ : SRMux
    port map (
            O => \N__27074\,
            I => \N__26920\
        );

    \I__6454\ : SRMux
    port map (
            O => \N__27073\,
            I => \N__26920\
        );

    \I__6453\ : SRMux
    port map (
            O => \N__27072\,
            I => \N__26920\
        );

    \I__6452\ : SRMux
    port map (
            O => \N__27071\,
            I => \N__26920\
        );

    \I__6451\ : SRMux
    port map (
            O => \N__27070\,
            I => \N__26920\
        );

    \I__6450\ : SRMux
    port map (
            O => \N__27069\,
            I => \N__26920\
        );

    \I__6449\ : SRMux
    port map (
            O => \N__27068\,
            I => \N__26920\
        );

    \I__6448\ : SRMux
    port map (
            O => \N__27067\,
            I => \N__26920\
        );

    \I__6447\ : SRMux
    port map (
            O => \N__27066\,
            I => \N__26920\
        );

    \I__6446\ : SRMux
    port map (
            O => \N__27065\,
            I => \N__26920\
        );

    \I__6445\ : SRMux
    port map (
            O => \N__27064\,
            I => \N__26920\
        );

    \I__6444\ : SRMux
    port map (
            O => \N__27063\,
            I => \N__26920\
        );

    \I__6443\ : GlobalMux
    port map (
            O => \N__26920\,
            I => \N__26917\
        );

    \I__6442\ : gio2CtrlBuf
    port map (
            O => \N__26917\,
            I => reset_n_i_g
        );

    \I__6441\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__26908\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_22\
        );

    \I__6438\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26901\
        );

    \I__6437\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26891\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__26901\,
            I => \N__26888\
        );

    \I__6435\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26873\
        );

    \I__6434\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26873\
        );

    \I__6433\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26873\
        );

    \I__6432\ : InMux
    port map (
            O => \N__26897\,
            I => \N__26873\
        );

    \I__6431\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26873\
        );

    \I__6430\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26873\
        );

    \I__6429\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26873\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26869\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__26888\,
            I => \N__26864\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__26873\,
            I => \N__26864\
        );

    \I__6425\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26855\
        );

    \I__6424\ : Span4Mux_s2_h
    port map (
            O => \N__26869\,
            I => \N__26850\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__26864\,
            I => \N__26850\
        );

    \I__6422\ : InMux
    port map (
            O => \N__26863\,
            I => \N__26837\
        );

    \I__6421\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26837\
        );

    \I__6420\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26837\
        );

    \I__6419\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26837\
        );

    \I__6418\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26837\
        );

    \I__6417\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26837\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__26855\,
            I => \ws2812.N_105\
        );

    \I__6415\ : Odrv4
    port map (
            O => \N__26850\,
            I => \ws2812.N_105\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__26837\,
            I => \ws2812.N_105\
        );

    \I__6413\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26827\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__26827\,
            I => \N__26824\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__26824\,
            I => rgb_data_out_23
        );

    \I__6410\ : CascadeMux
    port map (
            O => \N__26821\,
            I => \ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_\
        );

    \I__6409\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__26815\,
            I => \ws2812.N_117\
        );

    \I__6407\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26809\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__26809\,
            I => \N__26806\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__26806\,
            I => \N__26803\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__26803\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_3\
        );

    \I__6403\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__26797\,
            I => rgb_data_out_3
        );

    \I__6401\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26791\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26788\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__26788\,
            I => \N__26785\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__26785\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_19\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__26782\,
            I => \N__26779\
        );

    \I__6396\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26776\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__26776\,
            I => rgb_data_out_19
        );

    \I__6394\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26770\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__26770\,
            I => \N__26767\
        );

    \I__6392\ : Span12Mux_s4_h
    port map (
            O => \N__26767\,
            I => \N__26764\
        );

    \I__6391\ : Odrv12
    port map (
            O => \N__26764\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_7\
        );

    \I__6390\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__26758\,
            I => rgb_data_out_7
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__26755\,
            I => \N__26751\
        );

    \I__6387\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26746\
        );

    \I__6386\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26741\
        );

    \I__6385\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26736\
        );

    \I__6384\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26736\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26733\
        );

    \I__6382\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26728\
        );

    \I__6381\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26728\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__26741\,
            I => \ws2812.rgb_counter_4\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__26736\,
            I => \ws2812.rgb_counter_4\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__26733\,
            I => \ws2812.rgb_counter_4\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__26728\,
            I => \ws2812.rgb_counter_4\
        );

    \I__6376\ : CascadeMux
    port map (
            O => \N__26719\,
            I => \N__26716\
        );

    \I__6375\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26713\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26710\
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__26710\,
            I => rgb_data_out_22
        );

    \I__6372\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26704\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__26704\,
            I => \ws2812.rgb_data_pmux_6_i_m2_ns_1\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__26701\,
            I => \N__26698\
        );

    \I__6369\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26695\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__26695\,
            I => \ws2812.N_124\
        );

    \I__6367\ : InMux
    port map (
            O => \N__26692\,
            I => \ws2812.un1_rgb_counter_cry_3\
        );

    \I__6366\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26686\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__26686\,
            I => rgb_data_out_1
        );

    \I__6364\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26680\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__26680\,
            I => rgb_data_out_21
        );

    \I__6362\ : CascadeMux
    port map (
            O => \N__26677\,
            I => \ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_\
        );

    \I__6361\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__26671\,
            I => rgb_data_out_5
        );

    \I__6359\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__26662\,
            I => \ws2812.N_120\
        );

    \I__6356\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26656\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__26656\,
            I => \N__26653\
        );

    \I__6354\ : Span4Mux_s3_h
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__26650\,
            I => rgb_data_out_18
        );

    \I__6352\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__6350\ : Span4Mux_s2_h
    port map (
            O => \N__26641\,
            I => \N__26638\
        );

    \I__6349\ : Span4Mux_h
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__26635\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_2\
        );

    \I__6347\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__26629\,
            I => rgb_data_out_2
        );

    \I__6345\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26620\
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__26620\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_17\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__26617\,
            I => \N__26614\
        );

    \I__6341\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26611\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__26611\,
            I => rgb_data_out_17
        );

    \I__6339\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26605\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__26605\,
            I => \N__26602\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__26602\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_23\
        );

    \I__6336\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26596\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26593\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__26593\,
            I => \N__26590\
        );

    \I__6333\ : Odrv4
    port map (
            O => \N__26590\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_14\
        );

    \I__6332\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26581\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__26581\,
            I => rgb_data_out_14
        );

    \I__6329\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__26575\,
            I => \N__26572\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__26572\,
            I => \ws2812.data_RNOZ0Z_10\
        );

    \I__6326\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26566\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26563\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__26563\,
            I => \ws2812.data_RNOZ0Z_9\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__26560\,
            I => \N__26557\
        );

    \I__6322\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26554\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26551\
        );

    \I__6320\ : Odrv12
    port map (
            O => \N__26551\,
            I => \ws2812.data_RNOZ0Z_8\
        );

    \I__6319\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__26545\,
            I => \ws2812.N_135\
        );

    \I__6317\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__26539\,
            I => \ws2812.data_RNOZ0Z_2\
        );

    \I__6315\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_\
        );

    \I__6314\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26530\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__26530\,
            I => \ws2812.N_115\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__26527\,
            I => \N__26524\
        );

    \I__6311\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26521\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__26521\,
            I => \N__26518\
        );

    \I__6309\ : Odrv12
    port map (
            O => \N__26518\,
            I => rgb_data_out_16
        );

    \I__6308\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26512\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__26512\,
            I => \N__26509\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__26509\,
            I => rgb_data_out_0
        );

    \I__6305\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26500\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__26500\,
            I => rgb_data_out_20
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__26497\,
            I => \ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_\
        );

    \I__6301\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26491\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__26491\,
            I => \N__26488\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__26488\,
            I => rgb_data_out_4
        );

    \I__6298\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26482\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__26482\,
            I => \ws2812.N_127\
        );

    \I__6296\ : InMux
    port map (
            O => \N__26479\,
            I => \ws2812.un1_rgb_counter_cry_0\
        );

    \I__6295\ : InMux
    port map (
            O => \N__26476\,
            I => \ws2812.un1_rgb_counter_cry_1\
        );

    \I__6294\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__26467\,
            I => \N__26464\
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__26464\,
            I => \ws2812.rgb_counter_RNO_0Z0Z_3\
        );

    \I__6290\ : InMux
    port map (
            O => \N__26461\,
            I => \ws2812.un1_rgb_counter_cry_2\
        );

    \I__6289\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26455\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__26455\,
            I => \ws2812.un6_data_axb_8\
        );

    \I__6287\ : InMux
    port map (
            O => \N__26452\,
            I => \bfn_12_6_0_\
        );

    \I__6286\ : InMux
    port map (
            O => \N__26449\,
            I => \ws2812.un6_data_cry_8\
        );

    \I__6285\ : InMux
    port map (
            O => \N__26446\,
            I => \ws2812.un6_data_cry_9\
        );

    \I__6284\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26440\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__26437\,
            I => \ws2812.un6_data_axb_11\
        );

    \I__6281\ : InMux
    port map (
            O => \N__26434\,
            I => \ws2812.un6_data_cry_10\
        );

    \I__6280\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26428\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__26428\,
            I => \ws2812.data_RNOZ0Z_11\
        );

    \I__6278\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26422\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__26422\,
            I => \ws2812.data_RNOZ0Z_12\
        );

    \I__6276\ : CascadeMux
    port map (
            O => \N__26419\,
            I => \N__26416\
        );

    \I__6275\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26413\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__26413\,
            I => \ws2812.data_RNOZ0Z_13\
        );

    \I__6273\ : InMux
    port map (
            O => \N__26410\,
            I => \ws2812.un6_data_cry_11\
        );

    \I__6272\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26399\
        );

    \I__6270\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26396\
        );

    \I__6269\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26393\
        );

    \I__6268\ : Span4Mux_v
    port map (
            O => \N__26399\,
            I => \N__26389\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26384\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__26393\,
            I => \N__26384\
        );

    \I__6265\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26381\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__26389\,
            I => \ws2812.bit_counter_10\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__26384\,
            I => \ws2812.bit_counter_10\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__26381\,
            I => \ws2812.bit_counter_10\
        );

    \I__6261\ : InMux
    port map (
            O => \N__26374\,
            I => \N__26371\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__26371\,
            I => \ws2812.un6_data_axb_10\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__26368\,
            I => \N__26365\
        );

    \I__6258\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26361\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26355\
        );

    \I__6255\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26350\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__26355\,
            I => \N__26347\
        );

    \I__6253\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26344\
        );

    \I__6252\ : InMux
    port map (
            O => \N__26353\,
            I => \N__26341\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__26350\,
            I => \N__26338\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__26347\,
            I => \ws2812.bit_counter_9\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__26344\,
            I => \ws2812.bit_counter_9\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__26341\,
            I => \ws2812.bit_counter_9\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__26338\,
            I => \ws2812.bit_counter_9\
        );

    \I__6246\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__26326\,
            I => \ws2812.un6_data_axb_9\
        );

    \I__6244\ : InMux
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__26320\,
            I => \ws2812.data_RNOZ0Z_6\
        );

    \I__6242\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26314\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__26314\,
            I => \ws2812.data_RNOZ0Z_5\
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \N__26308\
        );

    \I__6239\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26305\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__26305\,
            I => \ws2812.data_5_iv_0_47_a2_0_a2_0\
        );

    \I__6237\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26299\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__26299\,
            I => \ws2812.data_5_iv_0_47_a2_0_a2_6_1\
        );

    \I__6235\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26293\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__26293\,
            I => \ws2812.data_5_iv_0_47_a2_0_a2_6\
        );

    \I__6233\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26286\
        );

    \I__6232\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26283\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__26286\,
            I => \ws2812.bit_counter_i_0\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__26283\,
            I => \ws2812.bit_counter_i_0\
        );

    \I__6229\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__26275\,
            I => \ws2812.un6_data_axb_1\
        );

    \I__6227\ : InMux
    port map (
            O => \N__26272\,
            I => \ws2812.un6_data_cry_0\
        );

    \I__6226\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__26266\,
            I => \ws2812.bit_counter_0_RNIQAT2Z0Z_0\
        );

    \I__6224\ : InMux
    port map (
            O => \N__26263\,
            I => \ws2812.un6_data_cry_1\
        );

    \I__6223\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__26257\,
            I => \ws2812.bit_counter_0_RNIRBT2Z0Z_1\
        );

    \I__6221\ : InMux
    port map (
            O => \N__26254\,
            I => \ws2812.un6_data_cry_2\
        );

    \I__6220\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__26248\,
            I => \N__26245\
        );

    \I__6218\ : Odrv4
    port map (
            O => \N__26245\,
            I => \ws2812.bit_counter_0_RNISCT2Z0Z_2\
        );

    \I__6217\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26236\
        );

    \I__6216\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26236\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__26236\,
            I => \N__26233\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__26233\,
            I => \ws2812.un6_data_cry_3_c_RNIKNFBZ0\
        );

    \I__6213\ : InMux
    port map (
            O => \N__26230\,
            I => \ws2812.un6_data_cry_3\
        );

    \I__6212\ : InMux
    port map (
            O => \N__26227\,
            I => \N__26224\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__26221\,
            I => \ws2812.bit_counter_0_RNITDT2Z0Z_3\
        );

    \I__6209\ : SRMux
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__26215\,
            I => \N__26204\
        );

    \I__6207\ : SRMux
    port map (
            O => \N__26214\,
            I => \N__26201\
        );

    \I__6206\ : SRMux
    port map (
            O => \N__26213\,
            I => \N__26198\
        );

    \I__6205\ : SRMux
    port map (
            O => \N__26212\,
            I => \N__26192\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__26211\,
            I => \N__26188\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__26210\,
            I => \N__26185\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__26209\,
            I => \N__26182\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__26208\,
            I => \N__26179\
        );

    \I__6200\ : SRMux
    port map (
            O => \N__26207\,
            I => \N__26174\
        );

    \I__6199\ : Span4Mux_s2_v
    port map (
            O => \N__26204\,
            I => \N__26163\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26163\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26163\
        );

    \I__6196\ : SRMux
    port map (
            O => \N__26197\,
            I => \N__26160\
        );

    \I__6195\ : SRMux
    port map (
            O => \N__26196\,
            I => \N__26157\
        );

    \I__6194\ : SRMux
    port map (
            O => \N__26195\,
            I => \N__26150\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__26192\,
            I => \N__26145\
        );

    \I__6192\ : SRMux
    port map (
            O => \N__26191\,
            I => \N__26142\
        );

    \I__6191\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26137\
        );

    \I__6190\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26137\
        );

    \I__6189\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26132\
        );

    \I__6188\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26132\
        );

    \I__6187\ : SRMux
    port map (
            O => \N__26178\,
            I => \N__26129\
        );

    \I__6186\ : SRMux
    port map (
            O => \N__26177\,
            I => \N__26126\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__26174\,
            I => \N__26120\
        );

    \I__6184\ : SRMux
    port map (
            O => \N__26173\,
            I => \N__26117\
        );

    \I__6183\ : SRMux
    port map (
            O => \N__26172\,
            I => \N__26114\
        );

    \I__6182\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26111\
        );

    \I__6181\ : SRMux
    port map (
            O => \N__26170\,
            I => \N__26108\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__26163\,
            I => \N__26101\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26101\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26101\
        );

    \I__6177\ : SRMux
    port map (
            O => \N__26156\,
            I => \N__26098\
        );

    \I__6176\ : SRMux
    port map (
            O => \N__26155\,
            I => \N__26094\
        );

    \I__6175\ : SRMux
    port map (
            O => \N__26154\,
            I => \N__26091\
        );

    \I__6174\ : SRMux
    port map (
            O => \N__26153\,
            I => \N__26088\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__26150\,
            I => \N__26085\
        );

    \I__6172\ : SRMux
    port map (
            O => \N__26149\,
            I => \N__26082\
        );

    \I__6171\ : SRMux
    port map (
            O => \N__26148\,
            I => \N__26079\
        );

    \I__6170\ : Span4Mux_v
    port map (
            O => \N__26145\,
            I => \N__26073\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__26142\,
            I => \N__26073\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__26137\,
            I => \N__26070\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26067\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26061\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26061\
        );

    \I__6164\ : SRMux
    port map (
            O => \N__26125\,
            I => \N__26058\
        );

    \I__6163\ : DummyBuf
    port map (
            O => \N__26124\,
            I => \N__26055\
        );

    \I__6162\ : DummyBuf
    port map (
            O => \N__26123\,
            I => \N__26052\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__26120\,
            I => \N__26045\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__26117\,
            I => \N__26045\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__26114\,
            I => \N__26045\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26040\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26040\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__26101\,
            I => \N__26035\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__26098\,
            I => \N__26035\
        );

    \I__6154\ : SRMux
    port map (
            O => \N__26097\,
            I => \N__26031\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26094\,
            I => \N__26028\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__26091\,
            I => \N__26023\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26023\
        );

    \I__6150\ : Span4Mux_s1_v
    port map (
            O => \N__26085\,
            I => \N__26016\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__26082\,
            I => \N__26016\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__26079\,
            I => \N__26016\
        );

    \I__6147\ : SRMux
    port map (
            O => \N__26078\,
            I => \N__26013\
        );

    \I__6146\ : Span4Mux_v
    port map (
            O => \N__26073\,
            I => \N__26006\
        );

    \I__6145\ : Span4Mux_s3_h
    port map (
            O => \N__26070\,
            I => \N__26006\
        );

    \I__6144\ : Span4Mux_s3_h
    port map (
            O => \N__26067\,
            I => \N__26006\
        );

    \I__6143\ : SRMux
    port map (
            O => \N__26066\,
            I => \N__26003\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__26061\,
            I => \N__25998\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__25998\
        );

    \I__6140\ : InMux
    port map (
            O => \N__26055\,
            I => \N__25995\
        );

    \I__6139\ : InMux
    port map (
            O => \N__26052\,
            I => \N__25992\
        );

    \I__6138\ : Span4Mux_v
    port map (
            O => \N__26045\,
            I => \N__25985\
        );

    \I__6137\ : Span4Mux_s3_h
    port map (
            O => \N__26040\,
            I => \N__25985\
        );

    \I__6136\ : Span4Mux_s3_v
    port map (
            O => \N__26035\,
            I => \N__25985\
        );

    \I__6135\ : SRMux
    port map (
            O => \N__26034\,
            I => \N__25982\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__26031\,
            I => \N__25979\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__26028\,
            I => \N__25976\
        );

    \I__6132\ : Span4Mux_v
    port map (
            O => \N__26023\,
            I => \N__25969\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__26016\,
            I => \N__25969\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__26013\,
            I => \N__25969\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__26006\,
            I => \N__25964\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__26003\,
            I => \N__25964\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__25998\,
            I => \N__25957\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__25995\,
            I => \N__25957\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25957\
        );

    \I__6124\ : Span4Mux_h
    port map (
            O => \N__25985\,
            I => \N__25952\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__25982\,
            I => \N__25952\
        );

    \I__6122\ : Sp12to4
    port map (
            O => \N__25979\,
            I => \N__25946\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25941\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__25969\,
            I => \N__25941\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__25964\,
            I => \N__25938\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__25957\,
            I => \N__25935\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__25952\,
            I => \N__25932\
        );

    \I__6116\ : SRMux
    port map (
            O => \N__25951\,
            I => \N__25929\
        );

    \I__6115\ : SRMux
    port map (
            O => \N__25950\,
            I => \N__25926\
        );

    \I__6114\ : SRMux
    port map (
            O => \N__25949\,
            I => \N__25923\
        );

    \I__6113\ : Odrv12
    port map (
            O => \N__25946\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6112\ : Odrv4
    port map (
            O => \N__25941\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__25938\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__25935\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__25932\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__25929\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__25926\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__25923\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25902\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__25905\,
            I => \N__25899\
        );

    \I__6103\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25894\
        );

    \I__6102\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25894\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__25894\,
            I => \N__25891\
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__25891\,
            I => \ws2812.un6_data_cry_4_c_RNIMQGBZ0\
        );

    \I__6099\ : InMux
    port map (
            O => \N__25888\,
            I => \ws2812.un6_data_cry_4\
        );

    \I__6098\ : InMux
    port map (
            O => \N__25885\,
            I => \N__25882\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__25882\,
            I => \ws2812.un6_data_axb_6\
        );

    \I__6096\ : InMux
    port map (
            O => \N__25879\,
            I => \ws2812.un6_data_cry_5\
        );

    \I__6095\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25873\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__25873\,
            I => \ws2812.un6_data_axb_7\
        );

    \I__6093\ : InMux
    port map (
            O => \N__25870\,
            I => \ws2812.un6_data_cry_6\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__25867\,
            I => \N__25863\
        );

    \I__6091\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25856\
        );

    \I__6090\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25845\
        );

    \I__6089\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25838\
        );

    \I__6088\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25838\
        );

    \I__6087\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25838\
        );

    \I__6086\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25833\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__25856\,
            I => \N__25830\
        );

    \I__6084\ : InMux
    port map (
            O => \N__25855\,
            I => \N__25821\
        );

    \I__6083\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25821\
        );

    \I__6082\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25821\
        );

    \I__6081\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25821\
        );

    \I__6080\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25816\
        );

    \I__6079\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25816\
        );

    \I__6078\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25811\
        );

    \I__6077\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25811\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__25845\,
            I => \N__25808\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25805\
        );

    \I__6074\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25802\
        );

    \I__6073\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25799\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__25833\,
            I => \N__25792\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__25830\,
            I => \N__25792\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25792\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25789\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__25811\,
            I => \N__25782\
        );

    \I__6067\ : Span4Mux_v
    port map (
            O => \N__25808\,
            I => \N__25782\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__25805\,
            I => \N__25782\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25777\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25777\
        );

    \I__6063\ : Span4Mux_h
    port map (
            O => \N__25792\,
            I => \N__25774\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__25789\,
            I => \demux.N_424_i_0_o2Z0Z_0\
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__25782\,
            I => \demux.N_424_i_0_o2Z0Z_0\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__25777\,
            I => \demux.N_424_i_0_o2Z0Z_0\
        );

    \I__6059\ : Odrv4
    port map (
            O => \N__25774\,
            I => \demux.N_424_i_0_o2Z0Z_0\
        );

    \I__6058\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25761\
        );

    \I__6057\ : InMux
    port map (
            O => \N__25764\,
            I => \N__25758\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25754\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25751\
        );

    \I__6054\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25748\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__25754\,
            I => \N__25744\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__25751\,
            I => \N__25739\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25739\
        );

    \I__6050\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25736\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__25744\,
            I => \N__25733\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__25739\,
            I => \N__25728\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25728\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__25733\,
            I => \demux.N_419_i_0_o2Z0Z_9\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__25728\,
            I => \demux.N_419_i_0_o2Z0Z_9\
        );

    \I__6044\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25719\
        );

    \I__6043\ : CascadeMux
    port map (
            O => \N__25722\,
            I => \N__25716\
        );

    \I__6042\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25712\
        );

    \I__6041\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25708\
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \N__25705\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25702\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__25711\,
            I => \N__25699\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__25708\,
            I => \N__25696\
        );

    \I__6036\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25693\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__25702\,
            I => \N__25690\
        );

    \I__6034\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25687\
        );

    \I__6033\ : Span4Mux_s3_h
    port map (
            O => \N__25696\,
            I => \N__25682\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__25693\,
            I => \N__25682\
        );

    \I__6031\ : Sp12to4
    port map (
            O => \N__25690\,
            I => \N__25677\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__25687\,
            I => \N__25677\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__25682\,
            I => \N__25674\
        );

    \I__6028\ : Span12Mux_v
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__6027\ : Sp12to4
    port map (
            O => \N__25674\,
            I => \N__25668\
        );

    \I__6026\ : Odrv12
    port map (
            O => \N__25671\,
            I => demux_data_in_5
        );

    \I__6025\ : Odrv12
    port map (
            O => \N__25668\,
            I => demux_data_in_5
        );

    \I__6024\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__6022\ : Span4Mux_s2_h
    port map (
            O => \N__25657\,
            I => \N__25651\
        );

    \I__6021\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25648\
        );

    \I__6020\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25645\
        );

    \I__6019\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25642\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__25651\,
            I => \demux.N_419_i_0_o2Z0Z_10\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__25648\,
            I => \demux.N_419_i_0_o2Z0Z_10\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__25645\,
            I => \demux.N_419_i_0_o2Z0Z_10\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__25642\,
            I => \demux.N_419_i_0_o2Z0Z_10\
        );

    \I__6014\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__25627\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_5\
        );

    \I__6011\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25619\
        );

    \I__6010\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25616\
        );

    \I__6009\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25613\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25610\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25607\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25604\
        );

    \I__6005\ : Span4Mux_s3_h
    port map (
            O => \N__25610\,
            I => \N__25600\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__25607\,
            I => \N__25597\
        );

    \I__6003\ : Span4Mux_s3_h
    port map (
            O => \N__25604\,
            I => \N__25594\
        );

    \I__6002\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25591\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__25600\,
            I => \demux.N_420_i_0_o2Z0Z_8\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__25597\,
            I => \demux.N_420_i_0_o2Z0Z_8\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__25594\,
            I => \demux.N_420_i_0_o2Z0Z_8\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__25591\,
            I => \demux.N_420_i_0_o2Z0Z_8\
        );

    \I__5997\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25578\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25575\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__25578\,
            I => \N__25571\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__25575\,
            I => \N__25567\
        );

    \I__5993\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25564\
        );

    \I__5992\ : Span4Mux_v
    port map (
            O => \N__25571\,
            I => \N__25561\
        );

    \I__5991\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25558\
        );

    \I__5990\ : Span4Mux_v
    port map (
            O => \N__25567\,
            I => \N__25553\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__25564\,
            I => \N__25553\
        );

    \I__5988\ : Sp12to4
    port map (
            O => \N__25561\,
            I => \N__25548\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__25558\,
            I => \N__25548\
        );

    \I__5986\ : Span4Mux_h
    port map (
            O => \N__25553\,
            I => \N__25545\
        );

    \I__5985\ : Odrv12
    port map (
            O => \N__25548\,
            I => \demux.N_420_i_0_o2Z0Z_9\
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__25545\,
            I => \demux.N_420_i_0_o2Z0Z_9\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__25540\,
            I => \N__25535\
        );

    \I__5982\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25531\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__25538\,
            I => \N__25528\
        );

    \I__5980\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25525\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__25534\,
            I => \N__25522\
        );

    \I__5978\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25519\
        );

    \I__5977\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25516\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__25525\,
            I => \N__25513\
        );

    \I__5975\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25510\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__25519\,
            I => \N__25507\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25504\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__25513\,
            I => \N__25499\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25499\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__25507\,
            I => \N__25494\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__25504\,
            I => \N__25494\
        );

    \I__5968\ : Span4Mux_h
    port map (
            O => \N__25499\,
            I => \N__25491\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__25494\,
            I => \demux.N_420_i_0_aZ0Z3\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__25491\,
            I => \demux.N_420_i_0_aZ0Z3\
        );

    \I__5965\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25481\
        );

    \I__5964\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25478\
        );

    \I__5963\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25474\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__25481\,
            I => \N__25471\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__25478\,
            I => \N__25468\
        );

    \I__5960\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25465\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__25474\,
            I => \N__25460\
        );

    \I__5958\ : Span4Mux_s3_h
    port map (
            O => \N__25471\,
            I => \N__25460\
        );

    \I__5957\ : Span4Mux_s3_h
    port map (
            O => \N__25468\,
            I => \N__25457\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__25465\,
            I => \demux.N_420_i_0_o2Z0Z_7\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__25460\,
            I => \demux.N_420_i_0_o2Z0Z_7\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__25457\,
            I => \demux.N_420_i_0_o2Z0Z_7\
        );

    \I__5953\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25444\
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__25444\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_4\
        );

    \I__5950\ : CEMux
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25434\
        );

    \I__5948\ : CEMux
    port map (
            O => \N__25437\,
            I => \N__25431\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__25434\,
            I => \N__25425\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25425\
        );

    \I__5945\ : CEMux
    port map (
            O => \N__25430\,
            I => \N__25422\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__25425\,
            I => \N__25417\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__25422\,
            I => \N__25417\
        );

    \I__5942\ : Span4Mux_h
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__25414\,
            I => \N__25411\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__25411\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1\
        );

    \I__5939\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25404\
        );

    \I__5938\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25390\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__25404\,
            I => \N__25387\
        );

    \I__5936\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25370\
        );

    \I__5935\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25370\
        );

    \I__5934\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25370\
        );

    \I__5933\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25370\
        );

    \I__5932\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25370\
        );

    \I__5931\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25370\
        );

    \I__5930\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25370\
        );

    \I__5929\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25370\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__25395\,
            I => \N__25366\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__25394\,
            I => \N__25362\
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__25393\,
            I => \N__25357\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25352\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__25387\,
            I => \N__25347\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__25370\,
            I => \N__25347\
        );

    \I__5922\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25342\
        );

    \I__5921\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25342\
        );

    \I__5920\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25339\
        );

    \I__5919\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25326\
        );

    \I__5918\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25326\
        );

    \I__5917\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25326\
        );

    \I__5916\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25326\
        );

    \I__5915\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25326\
        );

    \I__5914\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25326\
        );

    \I__5913\ : Span4Mux_v
    port map (
            O => \N__25352\,
            I => \N__25319\
        );

    \I__5912\ : Span4Mux_h
    port map (
            O => \N__25347\,
            I => \N__25319\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__25342\,
            I => \N__25319\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__25339\,
            I => \ws2812.stateZ0Z_1\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__25326\,
            I => \ws2812.stateZ0Z_1\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__25319\,
            I => \ws2812.stateZ0Z_1\
        );

    \I__5907\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25306\
        );

    \I__5906\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25306\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__25306\,
            I => \ws2812.state_ns_0_i_o2_8_0\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__25303\,
            I => \N__25300\
        );

    \I__5903\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__25297\,
            I => \N__25291\
        );

    \I__5901\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25288\
        );

    \I__5900\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25283\
        );

    \I__5899\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25283\
        );

    \I__5898\ : Odrv12
    port map (
            O => \N__25291\,
            I => \ws2812.bit_counterZ0Z_1\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__25288\,
            I => \ws2812.bit_counterZ0Z_1\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__25283\,
            I => \ws2812.bit_counterZ0Z_1\
        );

    \I__5895\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25271\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__25275\,
            I => \N__25267\
        );

    \I__5893\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25264\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25261\
        );

    \I__5891\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25258\
        );

    \I__5890\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25253\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__25264\,
            I => \N__25248\
        );

    \I__5888\ : Span4Mux_v
    port map (
            O => \N__25261\,
            I => \N__25248\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25245\
        );

    \I__5886\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25240\
        );

    \I__5885\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25240\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__25253\,
            I => \ws2812.bit_counterZ0Z_0\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__25248\,
            I => \ws2812.bit_counterZ0Z_0\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__25245\,
            I => \ws2812.bit_counterZ0Z_0\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__25240\,
            I => \ws2812.bit_counterZ0Z_0\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__25231\,
            I => \N__25227\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__25230\,
            I => \N__25223\
        );

    \I__5878\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25220\
        );

    \I__5877\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25215\
        );

    \I__5876\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25215\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__25220\,
            I => \N__25212\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__25215\,
            I => \N__25209\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__25212\,
            I => \ws2812.bit_counter_11\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__25209\,
            I => \ws2812.bit_counter_11\
        );

    \I__5871\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25201\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__25198\,
            I => \ws2812.bit_counter_0_RNO_0Z0Z_4\
        );

    \I__5868\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25192\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__25192\,
            I => \ws2812.bit_counter_0_RNO_0Z0Z_0\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__5865\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__25183\,
            I => \N__25177\
        );

    \I__5863\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25170\
        );

    \I__5862\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25170\
        );

    \I__5861\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25170\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__25177\,
            I => \ws2812.bit_counterZ0Z_2\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__25170\,
            I => \ws2812.bit_counterZ0Z_2\
        );

    \I__5858\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25162\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__25162\,
            I => \N__25159\
        );

    \I__5856\ : Span4Mux_v
    port map (
            O => \N__25159\,
            I => \N__25156\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__25156\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_13\
        );

    \I__5854\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25150\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__25150\,
            I => rgb_data_out_13
        );

    \I__5852\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25144\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__25138\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_11\
        );

    \I__5848\ : InMux
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__25129\,
            I => rgb_data_out_11
        );

    \I__5845\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25123\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__25123\,
            I => \N__25120\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__25117\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_9\
        );

    \I__5841\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25111\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__25111\,
            I => \N__25108\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__25108\,
            I => rgb_data_out_9
        );

    \I__5838\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25099\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__25099\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_1\
        );

    \I__5835\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25090\
        );

    \I__5833\ : Span4Mux_s3_h
    port map (
            O => \N__25090\,
            I => \N__25087\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__25087\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_21\
        );

    \I__5831\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__25081\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_20\
        );

    \I__5829\ : CEMux
    port map (
            O => \N__25078\,
            I => \N__25074\
        );

    \I__5828\ : CEMux
    port map (
            O => \N__25077\,
            I => \N__25071\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25068\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25065\
        );

    \I__5825\ : Span4Mux_s3_h
    port map (
            O => \N__25068\,
            I => \N__25062\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__25065\,
            I => \N__25059\
        );

    \I__5823\ : Span4Mux_v
    port map (
            O => \N__25062\,
            I => \N__25053\
        );

    \I__5822\ : Span4Mux_s3_h
    port map (
            O => \N__25059\,
            I => \N__25053\
        );

    \I__5821\ : CEMux
    port map (
            O => \N__25058\,
            I => \N__25050\
        );

    \I__5820\ : Span4Mux_h
    port map (
            O => \N__25053\,
            I => \N__25047\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__25050\,
            I => \N__25044\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__25047\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1\
        );

    \I__5817\ : Odrv12
    port map (
            O => \N__25044\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1\
        );

    \I__5816\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25036\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__25036\,
            I => \N__25033\
        );

    \I__5814\ : Span4Mux_s3_h
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__25030\,
            I => rgb_data_out_12
        );

    \I__5812\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25024\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__25024\,
            I => \N__25021\
        );

    \I__5810\ : Span4Mux_s3_h
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__25018\,
            I => rgb_data_out_15
        );

    \I__5808\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25012\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25009\
        );

    \I__5806\ : Span4Mux_s3_h
    port map (
            O => \N__25009\,
            I => \N__25006\
        );

    \I__5805\ : Odrv4
    port map (
            O => \N__25006\,
            I => rgb_data_out_10
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__25003\,
            I => \ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_\
        );

    \I__5803\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__24997\,
            I => \ws2812.rgb_counter_RNI2H7OZ0Z_2\
        );

    \I__5801\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__24991\,
            I => \ws2812.rgb_counter_RNIFI3MZ0Z_2\
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__24988\,
            I => \ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_\
        );

    \I__5798\ : CascadeMux
    port map (
            O => \N__24985\,
            I => \ws2812.N_108_cascade_\
        );

    \I__5797\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24976\
        );

    \I__5796\ : InMux
    port map (
            O => \N__24981\,
            I => \N__24976\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__24976\,
            I => \ws2812.N_107\
        );

    \I__5794\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24970\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__24970\,
            I => \ws2812.rgb_counter_RNI4J7OZ0Z_2\
        );

    \I__5792\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__5790\ : Span4Mux_h
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__24958\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_8\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__24952\,
            I => rgb_data_out_8
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \N__24946\
        );

    \I__5785\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__24940\,
            I => \ws2812.bit_counter_RNI9RQB3Z0Z_5\
        );

    \I__5782\ : InMux
    port map (
            O => \N__24937\,
            I => \ws2812.un1_bit_counter_12_cry_8\
        );

    \I__5781\ : CascadeMux
    port map (
            O => \N__24934\,
            I => \N__24931\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24925\
        );

    \I__5778\ : Odrv12
    port map (
            O => \N__24925\,
            I => \ws2812.bit_counter_0_RNING643Z0Z_4\
        );

    \I__5777\ : InMux
    port map (
            O => \N__24922\,
            I => \ws2812.un1_bit_counter_12_cry_9\
        );

    \I__5776\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24916\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__24913\,
            I => \ws2812.un1_bit_counter_12_axb_11\
        );

    \I__5773\ : InMux
    port map (
            O => \N__24910\,
            I => \ws2812.un1_bit_counter_12_cry_10\
        );

    \I__5772\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__5771\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24901\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__24901\,
            I => \N__24898\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__24898\,
            I => \ws2812.state_ns_0_i_o2_7_0\
        );

    \I__5768\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24890\
        );

    \I__5767\ : InMux
    port map (
            O => \N__24894\,
            I => \N__24884\
        );

    \I__5766\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24884\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24881\
        );

    \I__5764\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24878\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24875\
        );

    \I__5762\ : Odrv12
    port map (
            O => \N__24881\,
            I => \ws2812.bit_counterZ0Z_4\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__24878\,
            I => \ws2812.bit_counterZ0Z_4\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__24875\,
            I => \ws2812.bit_counterZ0Z_4\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__24868\,
            I => \N__24865\
        );

    \I__5758\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24860\
        );

    \I__5757\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24854\
        );

    \I__5756\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24854\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__24860\,
            I => \N__24851\
        );

    \I__5754\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24848\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24845\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__24851\,
            I => \ws2812.bit_counterZ0Z_5\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__24848\,
            I => \ws2812.bit_counterZ0Z_5\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__24845\,
            I => \ws2812.bit_counterZ0Z_5\
        );

    \I__5749\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24835\,
            I => \N__24829\
        );

    \I__5747\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24826\
        );

    \I__5746\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24821\
        );

    \I__5745\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24821\
        );

    \I__5744\ : Odrv12
    port map (
            O => \N__24829\,
            I => \ws2812.bit_counter_8\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__24826\,
            I => \ws2812.bit_counter_8\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__24821\,
            I => \ws2812.bit_counter_8\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__24814\,
            I => \ws2812.N_52_cascade_\
        );

    \I__5740\ : IoInMux
    port map (
            O => \N__24811\,
            I => \N__24808\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__24808\,
            I => \N__24805\
        );

    \I__5738\ : Span4Mux_s3_v
    port map (
            O => \N__24805\,
            I => \N__24801\
        );

    \I__5737\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24798\
        );

    \I__5736\ : Odrv4
    port map (
            O => \N__24801\,
            I => led
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__24798\,
            I => led
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__24793\,
            I => \N__24790\
        );

    \I__5733\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24784\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__24784\,
            I => \ws2812.bit_counter_RNI5NQB3Z0Z_1\
        );

    \I__5730\ : InMux
    port map (
            O => \N__24781\,
            I => \ws2812.un1_bit_counter_12_cry_0\
        );

    \I__5729\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24775\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__24775\,
            I => \ws2812.bit_counter_0_RNIJC643Z0Z_0\
        );

    \I__5727\ : InMux
    port map (
            O => \N__24772\,
            I => \ws2812.un1_bit_counter_12_cry_1\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__5725\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24761\
        );

    \I__5724\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24755\
        );

    \I__5723\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24755\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24752\
        );

    \I__5721\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24749\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24746\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__24752\,
            I => \N__24741\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24741\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__24746\,
            I => \N__24738\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__24741\,
            I => \ws2812.bit_counterZ0Z_3\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__24738\,
            I => \ws2812.bit_counterZ0Z_3\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__24733\,
            I => \N__24730\
        );

    \I__5713\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__24727\,
            I => \N__24724\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__24724\,
            I => \ws2812.bit_counter_0_RNIKD643Z0Z_1\
        );

    \I__5710\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24718\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__24718\,
            I => \N__24715\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__24715\,
            I => \ws2812.bit_counter_0_RNO_0Z0Z_1\
        );

    \I__5707\ : InMux
    port map (
            O => \N__24712\,
            I => \ws2812.un1_bit_counter_12_cry_2\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__24709\,
            I => \N__24706\
        );

    \I__5705\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__24703\,
            I => \N__24700\
        );

    \I__5703\ : Odrv4
    port map (
            O => \N__24700\,
            I => \ws2812.bit_counter_0_RNILE643Z0Z_2\
        );

    \I__5702\ : InMux
    port map (
            O => \N__24697\,
            I => \ws2812.un1_bit_counter_12_cry_3\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__5700\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24685\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__24685\,
            I => \ws2812.bit_counter_0_RNIMF643Z0Z_3\
        );

    \I__5697\ : InMux
    port map (
            O => \N__24682\,
            I => \ws2812.un1_bit_counter_12_cry_4\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__24679\,
            I => \N__24676\
        );

    \I__5695\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24673\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__5693\ : Span4Mux_h
    port map (
            O => \N__24670\,
            I => \N__24667\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__24667\,
            I => \ws2812.bit_counter_RNI6OQB3Z0Z_2\
        );

    \I__5691\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24661\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__24661\,
            I => \N__24658\
        );

    \I__5689\ : Span12Mux_s9_v
    port map (
            O => \N__24658\,
            I => \N__24652\
        );

    \I__5688\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24649\
        );

    \I__5687\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24644\
        );

    \I__5686\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24644\
        );

    \I__5685\ : Odrv12
    port map (
            O => \N__24652\,
            I => \ws2812.bit_counter_6\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__24649\,
            I => \ws2812.bit_counter_6\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__24644\,
            I => \ws2812.bit_counter_6\
        );

    \I__5682\ : InMux
    port map (
            O => \N__24637\,
            I => \ws2812.un1_bit_counter_12_cry_5\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__24634\,
            I => \N__24631\
        );

    \I__5680\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__5678\ : Span4Mux_s3_h
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__24622\,
            I => \ws2812.bit_counter_RNI7PQB3Z0Z_3\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__24619\,
            I => \N__24616\
        );

    \I__5675\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__24613\,
            I => \N__24609\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__24612\,
            I => \N__24604\
        );

    \I__5672\ : Span4Mux_v
    port map (
            O => \N__24609\,
            I => \N__24601\
        );

    \I__5671\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24598\
        );

    \I__5670\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24593\
        );

    \I__5669\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24593\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__24601\,
            I => \ws2812.bit_counter_7\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__24598\,
            I => \ws2812.bit_counter_7\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__24593\,
            I => \ws2812.bit_counter_7\
        );

    \I__5665\ : InMux
    port map (
            O => \N__24586\,
            I => \ws2812.un1_bit_counter_12_cry_6\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__5663\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24577\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__24574\,
            I => \ws2812.bit_counter_RNI8QQB3Z0Z_4\
        );

    \I__5660\ : InMux
    port map (
            O => \N__24571\,
            I => \bfn_11_6_0_\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__24568\,
            I => \ws2812.state_ns_0_i_o2_6_0_cascade_\
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__24565\,
            I => \ws2812.N_105_cascade_\
        );

    \I__5657\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__24559\,
            I => \ws2812.state_ns_0_i_o2_6_0\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__24556\,
            I => \N__24553\
        );

    \I__5654\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24550\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__24547\,
            I => \ws2812.un1_bit_counter_12_cry_0_c_RNOZ0\
        );

    \I__5651\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__24538\,
            I => \N__24535\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__24535\,
            I => demux_data_in_101
        );

    \I__5647\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__24529\,
            I => demux_data_in_21
        );

    \I__5645\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24523\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__24523\,
            I => \demux.N_419_i_0_o2Z0Z_4\
        );

    \I__5643\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__5641\ : Span4Mux_v
    port map (
            O => \N__24514\,
            I => \N__24511\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__24511\,
            I => demux_data_in_100
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24499\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__24507\,
            I => \N__24496\
        );

    \I__5637\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24493\
        );

    \I__5636\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24488\
        );

    \I__5635\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24488\
        );

    \I__5634\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24479\
        );

    \I__5633\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24479\
        );

    \I__5632\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24479\
        );

    \I__5631\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24479\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24475\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__24488\,
            I => \N__24472\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24469\
        );

    \I__5627\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24466\
        );

    \I__5626\ : Span4Mux_h
    port map (
            O => \N__24475\,
            I => \N__24463\
        );

    \I__5625\ : Span4Mux_h
    port map (
            O => \N__24472\,
            I => \N__24458\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__24469\,
            I => \N__24458\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__24466\,
            I => \demux.N_424_i_0_a2Z0Z_3\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__24463\,
            I => \demux.N_424_i_0_a2Z0Z_3\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__24458\,
            I => \demux.N_424_i_0_a2Z0Z_3\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__5619\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24445\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__24445\,
            I => \N__24442\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__24439\,
            I => demux_data_in_20
        );

    \I__5615\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24427\
        );

    \I__5614\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24424\
        );

    \I__5613\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24421\
        );

    \I__5612\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24412\
        );

    \I__5611\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24412\
        );

    \I__5610\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24412\
        );

    \I__5609\ : InMux
    port map (
            O => \N__24430\,
            I => \N__24412\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24408\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__24424\,
            I => \N__24405\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24402\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24399\
        );

    \I__5604\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24396\
        );

    \I__5603\ : Span4Mux_h
    port map (
            O => \N__24408\,
            I => \N__24393\
        );

    \I__5602\ : Span4Mux_h
    port map (
            O => \N__24405\,
            I => \N__24390\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__24402\,
            I => \N__24385\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__24399\,
            I => \N__24385\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__24396\,
            I => \demux.N_424_i_0_a2Z0Z_10\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__24393\,
            I => \demux.N_424_i_0_a2Z0Z_10\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__24390\,
            I => \demux.N_424_i_0_a2Z0Z_10\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__24385\,
            I => \demux.N_424_i_0_a2Z0Z_10\
        );

    \I__5595\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24373\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__24370\,
            I => \N__24367\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__5591\ : Odrv4
    port map (
            O => \N__24364\,
            I => demux_data_in_68
        );

    \I__5590\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24355\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__24360\,
            I => \N__24350\
        );

    \I__5588\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24344\
        );

    \I__5587\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24344\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24341\
        );

    \I__5585\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24338\
        );

    \I__5584\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24335\
        );

    \I__5583\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24330\
        );

    \I__5582\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24330\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__24344\,
            I => \N__24327\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__24341\,
            I => \N__24321\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24321\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24318\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24315\
        );

    \I__5576\ : Span4Mux_s3_v
    port map (
            O => \N__24327\,
            I => \N__24312\
        );

    \I__5575\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24309\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__24321\,
            I => \N__24304\
        );

    \I__5573\ : Span4Mux_s3_v
    port map (
            O => \N__24318\,
            I => \N__24304\
        );

    \I__5572\ : Span4Mux_h
    port map (
            O => \N__24315\,
            I => \N__24301\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__24312\,
            I => \demux.N_424_i_0_a2Z0Z_9\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__24309\,
            I => \demux.N_424_i_0_a2Z0Z_9\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__24304\,
            I => \demux.N_424_i_0_a2Z0Z_9\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__24301\,
            I => \demux.N_424_i_0_a2Z0Z_9\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__24292\,
            I => \demux.N_420_i_0_o2Z0Z_4_cascade_\
        );

    \I__5566\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__24280\,
            I => \demux.N_420_i_0_a3Z0Z_7\
        );

    \I__5562\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__5560\ : Span12Mux_s9_h
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__5559\ : Odrv12
    port map (
            O => \N__24268\,
            I => miso_data_in_5
        );

    \I__5558\ : InMux
    port map (
            O => \N__24265\,
            I => \N__24260\
        );

    \I__5557\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24257\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \N__24253\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24248\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24248\
        );

    \I__5553\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24245\
        );

    \I__5552\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24242\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__24248\,
            I => \N__24239\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24236\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24233\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__24239\,
            I => \N__24230\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__24236\,
            I => \N__24225\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__24233\,
            I => \N__24225\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__24230\,
            I => \demux.N_421_i_0_o2Z0Z_9\
        );

    \I__5544\ : Odrv4
    port map (
            O => \N__24225\,
            I => \demux.N_421_i_0_o2Z0Z_9\
        );

    \I__5543\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24215\
        );

    \I__5542\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24212\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__24218\,
            I => \N__24208\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24205\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__24212\,
            I => \N__24202\
        );

    \I__5538\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24199\
        );

    \I__5537\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24196\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__24205\,
            I => \N__24187\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__24202\,
            I => \N__24187\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__24199\,
            I => \N__24187\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24187\
        );

    \I__5532\ : Span4Mux_v
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__24184\,
            I => \N__24181\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__24181\,
            I => demux_data_in_3
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__24178\,
            I => \N__24173\
        );

    \I__5528\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24169\
        );

    \I__5527\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24166\
        );

    \I__5526\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24163\
        );

    \I__5525\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24160\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24157\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24152\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__24163\,
            I => \N__24152\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__24160\,
            I => \demux.N_421_i_0_o2Z0Z_10\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__24157\,
            I => \demux.N_421_i_0_o2Z0Z_10\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__24152\,
            I => \demux.N_421_i_0_o2Z0Z_10\
        );

    \I__5518\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24142\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__24142\,
            I => \N__24139\
        );

    \I__5516\ : Odrv12
    port map (
            O => \N__24139\,
            I => miso_data_in_3
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__24136\,
            I => \N__24132\
        );

    \I__5514\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24128\
        );

    \I__5513\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24125\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24122\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24118\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__24125\,
            I => \N__24113\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__24122\,
            I => \N__24113\
        );

    \I__5508\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24110\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__24118\,
            I => \N__24103\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__24113\,
            I => \N__24103\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24103\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__24100\,
            I => \demux.N_423_i_0_o2Z0Z_9\
        );

    \I__5502\ : CascadeMux
    port map (
            O => \N__24097\,
            I => \N__24094\
        );

    \I__5501\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24089\
        );

    \I__5500\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24086\
        );

    \I__5499\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24082\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24077\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__24086\,
            I => \N__24077\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__24085\,
            I => \N__24074\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24071\
        );

    \I__5494\ : Span4Mux_v
    port map (
            O => \N__24077\,
            I => \N__24068\
        );

    \I__5493\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24065\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__24071\,
            I => \N__24062\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__24068\,
            I => \N__24057\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__24065\,
            I => \N__24057\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__24062\,
            I => \N__24054\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__24057\,
            I => \N__24051\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__24054\,
            I => demux_data_in_1
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__24051\,
            I => demux_data_in_1
        );

    \I__5485\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24040\
        );

    \I__5484\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24037\
        );

    \I__5483\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24034\
        );

    \I__5482\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24031\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__24040\,
            I => \demux.N_423_i_0_o2Z0Z_10\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__24037\,
            I => \demux.N_423_i_0_o2Z0Z_10\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__24034\,
            I => \demux.N_423_i_0_o2Z0Z_10\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__24031\,
            I => \demux.N_423_i_0_o2Z0Z_10\
        );

    \I__5477\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24019\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__5475\ : Odrv12
    port map (
            O => \N__24016\,
            I => miso_data_in_1
        );

    \I__5474\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24010\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__24007\,
            I => \N__24004\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__24004\,
            I => \N__24001\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__24001\,
            I => miso_data_in_4
        );

    \I__5469\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__23995\,
            I => \N__23988\
        );

    \I__5467\ : CEMux
    port map (
            O => \N__23994\,
            I => \N__23977\
        );

    \I__5466\ : CEMux
    port map (
            O => \N__23993\,
            I => \N__23977\
        );

    \I__5465\ : CEMux
    port map (
            O => \N__23992\,
            I => \N__23977\
        );

    \I__5464\ : CEMux
    port map (
            O => \N__23991\,
            I => \N__23977\
        );

    \I__5463\ : Glb2LocalMux
    port map (
            O => \N__23988\,
            I => \N__23977\
        );

    \I__5462\ : GlobalMux
    port map (
            O => \N__23977\,
            I => \N__23974\
        );

    \I__5461\ : gio2CtrlBuf
    port map (
            O => \N__23974\,
            I => \sb_translator_1.state_g_1\
        );

    \I__5460\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23968\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__5458\ : Sp12to4
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__5457\ : Span12Mux_v
    port map (
            O => \N__23962\,
            I => \N__23959\
        );

    \I__5456\ : Odrv12
    port map (
            O => \N__23959\,
            I => demux_data_in_31
        );

    \I__5455\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23952\
        );

    \I__5454\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23946\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23943\
        );

    \I__5452\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23940\
        );

    \I__5451\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23935\
        );

    \I__5450\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23935\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__23946\,
            I => \N__23932\
        );

    \I__5448\ : Span4Mux_h
    port map (
            O => \N__23943\,
            I => \N__23923\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23923\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23923\
        );

    \I__5445\ : Span4Mux_h
    port map (
            O => \N__23932\,
            I => \N__23919\
        );

    \I__5444\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23914\
        );

    \I__5443\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23914\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__23923\,
            I => \N__23911\
        );

    \I__5441\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23908\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__23919\,
            I => \demux.N_424_i_0_a2Z0Z_1\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__23914\,
            I => \demux.N_424_i_0_a2Z0Z_1\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__23911\,
            I => \demux.N_424_i_0_a2Z0Z_1\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__23908\,
            I => \demux.N_424_i_0_a2Z0Z_1\
        );

    \I__5436\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23896\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23893\
        );

    \I__5434\ : Span12Mux_s10_h
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__5433\ : Odrv12
    port map (
            O => \N__23890\,
            I => demux_data_in_71
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__23887\,
            I => \demux.N_417_i_0_a3Z0Z_7_cascade_\
        );

    \I__5431\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23878\
        );

    \I__5430\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23875\
        );

    \I__5429\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23872\
        );

    \I__5428\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23869\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__23878\,
            I => \N__23860\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__23875\,
            I => \N__23860\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__23872\,
            I => \N__23860\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23860\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__23860\,
            I => \demux.N_417_i_0_o2Z0Z_8\
        );

    \I__5422\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23854\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__5420\ : Span4Mux_v
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__23848\,
            I => demux_data_in_103
        );

    \I__5418\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__23842\,
            I => demux_data_in_23
        );

    \I__5416\ : InMux
    port map (
            O => \N__23839\,
            I => \N__23836\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__23836\,
            I => \demux.N_417_i_0_o2Z0Z_4\
        );

    \I__5414\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__23827\,
            I => demux_data_in_18
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__23824\,
            I => \N__23821\
        );

    \I__5410\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23815\
        );

    \I__5408\ : Sp12to4
    port map (
            O => \N__23815\,
            I => \N__23812\
        );

    \I__5407\ : Odrv12
    port map (
            O => \N__23812\,
            I => demux_data_in_98
        );

    \I__5406\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__23800\,
            I => \demux.N_422_i_0_o2Z0Z_4\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__23797\,
            I => \demux.N_874_cascade_\
        );

    \I__5401\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23791\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__5397\ : Odrv4
    port map (
            O => \N__23782\,
            I => demux_data_in_4
        );

    \I__5396\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23775\
        );

    \I__5395\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23772\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__23775\,
            I => \N__23767\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23764\
        );

    \I__5392\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23761\
        );

    \I__5391\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23758\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__23767\,
            I => \N__23755\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__23764\,
            I => \N__23752\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__23761\,
            I => \N__23749\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__23758\,
            I => \N__23746\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__23755\,
            I => \N__23743\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__23752\,
            I => \N__23740\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__23749\,
            I => \N__23737\
        );

    \I__5383\ : Span4Mux_h
    port map (
            O => \N__23746\,
            I => \N__23734\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__23743\,
            I => \demux.N_417_i_0_o2Z0Z_9\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__23740\,
            I => \demux.N_417_i_0_o2Z0Z_9\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__23737\,
            I => \demux.N_417_i_0_o2Z0Z_9\
        );

    \I__5379\ : Odrv4
    port map (
            O => \N__23734\,
            I => \demux.N_417_i_0_o2Z0Z_9\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__23725\,
            I => \N__23722\
        );

    \I__5377\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23718\
        );

    \I__5376\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23715\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23709\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23709\
        );

    \I__5373\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23706\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__23709\,
            I => \demux.N_888\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__23706\,
            I => \demux.N_888\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__23701\,
            I => \N__23695\
        );

    \I__5369\ : CascadeMux
    port map (
            O => \N__23700\,
            I => \N__23692\
        );

    \I__5368\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23689\
        );

    \I__5367\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23686\
        );

    \I__5366\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23683\
        );

    \I__5365\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23680\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__23689\,
            I => \demux.N_417_i_0_o2Z0Z_7\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__23686\,
            I => \demux.N_417_i_0_o2Z0Z_7\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__23683\,
            I => \demux.N_417_i_0_o2Z0Z_7\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__23680\,
            I => \demux.N_417_i_0_o2Z0Z_7\
        );

    \I__5360\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__5358\ : Span12Mux_s5_h
    port map (
            O => \N__23665\,
            I => \N__23662\
        );

    \I__5357\ : Odrv12
    port map (
            O => \N__23662\,
            I => miso_data_in_7
        );

    \I__5356\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23655\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__23658\,
            I => \N__23652\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__23655\,
            I => \N__23649\
        );

    \I__5353\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23646\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__23649\,
            I => \N__23642\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23639\
        );

    \I__5350\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23636\
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__23642\,
            I => \demux.N_874\
        );

    \I__5348\ : Odrv12
    port map (
            O => \N__23639\,
            I => \demux.N_874\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__23636\,
            I => \demux.N_874\
        );

    \I__5346\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23622\
        );

    \I__5344\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23619\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__23622\,
            I => \N__23612\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__23619\,
            I => \N__23612\
        );

    \I__5341\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__5340\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23606\
        );

    \I__5339\ : Odrv4
    port map (
            O => \N__23612\,
            I => \demux.N_418_i_0_o2Z0Z_8\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__23609\,
            I => \demux.N_418_i_0_o2Z0Z_8\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__23606\,
            I => \demux.N_418_i_0_o2Z0Z_8\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__23599\,
            I => \N__23596\
        );

    \I__5335\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23592\
        );

    \I__5334\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__23592\,
            I => \N__23583\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__23589\,
            I => \N__23583\
        );

    \I__5331\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \N__23579\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__23583\,
            I => \N__23576\
        );

    \I__5329\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23573\
        );

    \I__5328\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23570\
        );

    \I__5327\ : Sp12to4
    port map (
            O => \N__23576\,
            I => \N__23563\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23563\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23563\
        );

    \I__5324\ : Odrv12
    port map (
            O => \N__23563\,
            I => \demux.N_418_i_0_o2Z0Z_9\
        );

    \I__5323\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23555\
        );

    \I__5322\ : InMux
    port map (
            O => \N__23559\,
            I => \N__23552\
        );

    \I__5321\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23548\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__23555\,
            I => \N__23543\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__23552\,
            I => \N__23543\
        );

    \I__5318\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23540\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__23548\,
            I => \demux.N_418_i_0_o2Z0Z_7\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__23543\,
            I => \demux.N_418_i_0_o2Z0Z_7\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__23540\,
            I => \demux.N_418_i_0_o2Z0Z_7\
        );

    \I__5314\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23530\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__5312\ : Odrv12
    port map (
            O => \N__23527\,
            I => miso_data_in_6
        );

    \I__5311\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23521\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__23521\,
            I => \N__23518\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__23518\,
            I => \N__23515\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__23515\,
            I => demux_data_in_14
        );

    \I__5307\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__23509\,
            I => \demux.N_880\
        );

    \I__5305\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23503\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__23500\,
            I => \N__23497\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__23497\,
            I => \N__23494\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__23491\,
            I => demux_data_in_36
        );

    \I__5299\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23482\
        );

    \I__5298\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23482\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23474\
        );

    \I__5296\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23469\
        );

    \I__5295\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23469\
        );

    \I__5294\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23466\
        );

    \I__5293\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23461\
        );

    \I__5292\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23461\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__23474\,
            I => \N__23456\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23456\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__23466\,
            I => \N__23453\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__23461\,
            I => \N__23449\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__23456\,
            I => \N__23444\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__23453\,
            I => \N__23444\
        );

    \I__5285\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23441\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__23449\,
            I => \demux.N_424_i_0_a2Z0Z_4\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__23444\,
            I => \demux.N_424_i_0_a2Z0Z_4\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__23441\,
            I => \demux.N_424_i_0_a2Z0Z_4\
        );

    \I__5281\ : CascadeMux
    port map (
            O => \N__23434\,
            I => \N__23430\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__23433\,
            I => \N__23427\
        );

    \I__5279\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23419\
        );

    \I__5278\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23419\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__23426\,
            I => \N__23416\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__23425\,
            I => \N__23413\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__23424\,
            I => \N__23409\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23405\
        );

    \I__5273\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23400\
        );

    \I__5272\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23400\
        );

    \I__5271\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23397\
        );

    \I__5270\ : InMux
    port map (
            O => \N__23409\,
            I => \N__23392\
        );

    \I__5269\ : InMux
    port map (
            O => \N__23408\,
            I => \N__23392\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__23405\,
            I => \N__23387\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__23400\,
            I => \N__23387\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__23397\,
            I => \N__23384\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__23392\,
            I => \demux.N_424_i_0_a2Z0Z_5\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__23387\,
            I => \demux.N_424_i_0_a2Z0Z_5\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__23384\,
            I => \demux.N_424_i_0_a2Z0Z_5\
        );

    \I__5262\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23374\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__23374\,
            I => demux_data_in_108
        );

    \I__5260\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23362\
        );

    \I__5259\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23357\
        );

    \I__5258\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23357\
        );

    \I__5257\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23352\
        );

    \I__5256\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23352\
        );

    \I__5255\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23347\
        );

    \I__5254\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23347\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23343\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__23357\,
            I => \N__23340\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__23352\,
            I => \N__23335\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__23347\,
            I => \N__23335\
        );

    \I__5249\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23332\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__23343\,
            I => \N__23327\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__23340\,
            I => \N__23327\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__23335\,
            I => \N__23324\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__23332\,
            I => \demux.N_424_i_0_a2Z0Z_11\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__23327\,
            I => \demux.N_424_i_0_a2Z0Z_11\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__23324\,
            I => \demux.N_424_i_0_a2Z0Z_11\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__23317\,
            I => \demux.N_420_i_0_o2Z0Z_0_cascade_\
        );

    \I__5241\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23311\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23308\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__23305\,
            I => demux_data_in_92
        );

    \I__5237\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23290\
        );

    \I__5235\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23287\
        );

    \I__5234\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23284\
        );

    \I__5233\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23281\
        );

    \I__5232\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23278\
        );

    \I__5231\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23273\
        );

    \I__5230\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23273\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__23290\,
            I => \N__23267\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23267\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__23284\,
            I => \N__23264\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23257\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__23278\,
            I => \N__23257\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23257\
        );

    \I__5223\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23254\
        );

    \I__5222\ : Span4Mux_v
    port map (
            O => \N__23267\,
            I => \N__23251\
        );

    \I__5221\ : Span4Mux_h
    port map (
            O => \N__23264\,
            I => \N__23248\
        );

    \I__5220\ : Span4Mux_v
    port map (
            O => \N__23257\,
            I => \N__23243\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23243\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__23251\,
            I => \demux.N_424_i_0_a2Z0Z_2\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__23248\,
            I => \demux.N_424_i_0_a2Z0Z_2\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__23243\,
            I => \demux.N_424_i_0_a2Z0Z_2\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__23230\,
            I => \N__23227\
        );

    \I__5212\ : Span4Mux_s3_h
    port map (
            O => \N__23227\,
            I => \N__23224\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__23224\,
            I => demux_data_in_12
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__23221\,
            I => \demux.N_420_i_0_o2Z0Z_1_cascade_\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23215\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__23212\,
            I => \demux.N_420_i_0_a3Z0Z_4\
        );

    \I__5206\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__5204\ : Sp12to4
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__23200\,
            I => demux_data_in_7
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__23197\,
            I => \demux.N_888_cascade_\
        );

    \I__5201\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23191\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23188\
        );

    \I__5199\ : Sp12to4
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__5198\ : Odrv12
    port map (
            O => \N__23185\,
            I => demux_data_in_6
        );

    \I__5197\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23179\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__23176\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_0\
        );

    \I__5194\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23170\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__23167\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_10\
        );

    \I__5191\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23161\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__23158\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_12\
        );

    \I__5188\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__23149\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_18\
        );

    \I__5185\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23143\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__23137\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_15\
        );

    \I__5181\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23131\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__23128\,
            I => \sb_translator_1.rgb_data_tmpZ0Z_16\
        );

    \I__5178\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__23119\,
            I => demux_data_in_94
        );

    \I__5175\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23113\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__23113\,
            I => demux_data_in_110
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__23110\,
            I => \demux.N_418_i_0_o2Z0Z_0_cascade_\
        );

    \I__5172\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23104\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__5168\ : Span4Mux_v
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__23092\,
            I => demux_data_in_38
        );

    \I__5166\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__5164\ : Span12Mux_s10_h
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__5163\ : Odrv12
    port map (
            O => \N__23080\,
            I => demux_data_in_46
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__23077\,
            I => \demux.N_418_i_0_o2Z0Z_1_cascade_\
        );

    \I__5161\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23068\
        );

    \I__5160\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23065\
        );

    \I__5159\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23061\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23058\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23050\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23050\
        );

    \I__5155\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23047\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23042\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23042\
        );

    \I__5152\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23037\
        );

    \I__5151\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23037\
        );

    \I__5150\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23034\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__23050\,
            I => \N__23031\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23028\
        );

    \I__5147\ : Span4Mux_v
    port map (
            O => \N__23042\,
            I => \N__23023\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23023\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__23034\,
            I => \N__23020\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__23031\,
            I => \demux.N_424_i_0_a2Z0Z_8\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__23028\,
            I => \demux.N_424_i_0_a2Z0Z_8\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__23023\,
            I => \demux.N_424_i_0_a2Z0Z_8\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__23020\,
            I => \demux.N_424_i_0_a2Z0Z_8\
        );

    \I__5140\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23005\
        );

    \I__5139\ : InMux
    port map (
            O => \N__23010\,
            I => \N__23000\
        );

    \I__5138\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23000\
        );

    \I__5137\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22994\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__23005\,
            I => \N__22991\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22988\
        );

    \I__5134\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22981\
        );

    \I__5133\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22981\
        );

    \I__5132\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22981\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__22994\,
            I => \N__22975\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__22991\,
            I => \N__22972\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__22988\,
            I => \N__22969\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__22981\,
            I => \N__22966\
        );

    \I__5127\ : InMux
    port map (
            O => \N__22980\,
            I => \N__22959\
        );

    \I__5126\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22959\
        );

    \I__5125\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22959\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__22975\,
            I => \N__22954\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__22972\,
            I => \N__22954\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__22969\,
            I => \sb_translator_1.stateZ0Z_6\
        );

    \I__5121\ : Odrv12
    port map (
            O => \N__22966\,
            I => \sb_translator_1.stateZ0Z_6\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__22959\,
            I => \sb_translator_1.stateZ0Z_6\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__22954\,
            I => \sb_translator_1.stateZ0Z_6\
        );

    \I__5118\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22941\
        );

    \I__5117\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22938\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22933\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22933\
        );

    \I__5114\ : Span4Mux_v
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__22930\,
            I => mosi_data_out_15
        );

    \I__5112\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22923\
        );

    \I__5111\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22920\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22916\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__22920\,
            I => \N__22913\
        );

    \I__5108\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22910\
        );

    \I__5107\ : Span4Mux_s2_h
    port map (
            O => \N__22916\,
            I => \N__22907\
        );

    \I__5106\ : Odrv12
    port map (
            O => \N__22913\,
            I => \sb_translator_1.cntZ0Z_7\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__22910\,
            I => \sb_translator_1.cntZ0Z_7\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__22907\,
            I => \sb_translator_1.cntZ0Z_7\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__5102\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__22891\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_7\
        );

    \I__5099\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__22879\,
            I => \ws2812.new_data_req_e_1\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \ws2812.N_140_cascade_\
        );

    \I__5094\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22870\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__22870\,
            I => \N__22866\
        );

    \I__5092\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__5091\ : Span12Mux_s8_v
    port map (
            O => \N__22866\,
            I => \N__22860\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__22863\,
            I => ws2812_next_led
        );

    \I__5089\ : Odrv12
    port map (
            O => \N__22860\,
            I => ws2812_next_led
        );

    \I__5088\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__22852\,
            I => \sb_translator_1.state56_a_5_8\
        );

    \I__5086\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22846\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__22846\,
            I => \sb_translator_1.state56_a_5_9\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__22843\,
            I => \sb_translator_1.N_318_i_i_o2_11_cascade_\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22837\,
            I => \sb_translator_1.state56_a_5_15\
        );

    \I__5081\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__22831\,
            I => \sb_translator_1.N_318_i_i_o2_14\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__5078\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22822\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__22822\,
            I => \N__22817\
        );

    \I__5076\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22812\
        );

    \I__5075\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22812\
        );

    \I__5074\ : Span4Mux_s3_v
    port map (
            O => \N__22817\,
            I => \N__22807\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22807\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__22804\,
            I => \N__22801\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__22801\,
            I => \sb_translator_1.state_RNII30CZ0Z_0\
        );

    \I__5069\ : IoInMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__22792\,
            I => \sb_translator_1.stateZ0Z_1\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__22789\,
            I => \N__22776\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__22788\,
            I => \N__22773\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__22787\,
            I => \N__22770\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__22786\,
            I => \N__22767\
        );

    \I__5062\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22756\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__22784\,
            I => \N__22753\
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22748\
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__22782\,
            I => \N__22745\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__22781\,
            I => \N__22742\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__22780\,
            I => \N__22739\
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__22779\,
            I => \N__22736\
        );

    \I__5055\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22725\
        );

    \I__5054\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22725\
        );

    \I__5053\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22725\
        );

    \I__5052\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22725\
        );

    \I__5051\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22716\
        );

    \I__5050\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22716\
        );

    \I__5049\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22716\
        );

    \I__5048\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22716\
        );

    \I__5047\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22713\
        );

    \I__5046\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22706\
        );

    \I__5045\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22706\
        );

    \I__5044\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22706\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22703\
        );

    \I__5042\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22696\
        );

    \I__5041\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22696\
        );

    \I__5040\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22696\
        );

    \I__5039\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22691\
        );

    \I__5038\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22691\
        );

    \I__5037\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22680\
        );

    \I__5036\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22680\
        );

    \I__5035\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22680\
        );

    \I__5034\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22680\
        );

    \I__5033\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22680\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22671\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22671\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22671\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__22706\,
            I => \N__22671\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__22703\,
            I => \N__22668\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22665\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22662\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22659\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__22671\,
            I => \N__22652\
        );

    \I__5023\ : Span4Mux_v
    port map (
            O => \N__22668\,
            I => \N__22652\
        );

    \I__5022\ : Span4Mux_h
    port map (
            O => \N__22665\,
            I => \N__22652\
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__22662\,
            I => mosi_data_out_23
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__22659\,
            I => mosi_data_out_23
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__22652\,
            I => mosi_data_out_23
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__22645\,
            I => \N__22640\
        );

    \I__5017\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22635\
        );

    \I__5016\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22632\
        );

    \I__5015\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22629\
        );

    \I__5014\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22624\
        );

    \I__5013\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22624\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22619\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__22632\,
            I => \N__22619\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__22629\,
            I => \N__22614\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22614\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__22619\,
            I => \N__22611\
        );

    \I__5007\ : Span12Mux_s9_h
    port map (
            O => \N__22614\,
            I => \N__22608\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__22611\,
            I => mosi_data_out_21
        );

    \I__5005\ : Odrv12
    port map (
            O => \N__22608\,
            I => mosi_data_out_21
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22599\
        );

    \I__5003\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22591\
        );

    \I__5002\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22591\
        );

    \I__5001\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22591\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__22591\,
            I => \N__22588\
        );

    \I__4999\ : Span12Mux_s9_h
    port map (
            O => \N__22588\,
            I => \N__22585\
        );

    \I__4998\ : Odrv12
    port map (
            O => \N__22585\,
            I => \sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0\
        );

    \I__4997\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__22579\,
            I => \N__22575\
        );

    \I__4995\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22572\
        );

    \I__4994\ : Span4Mux_h
    port map (
            O => \N__22575\,
            I => \N__22569\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__22572\,
            I => mosi_data_out_12
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__22569\,
            I => mosi_data_out_12
        );

    \I__4991\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22561\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22557\
        );

    \I__4989\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22553\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__22557\,
            I => \N__22550\
        );

    \I__4987\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22547\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22544\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__22550\,
            I => \sb_translator_1.cntZ0Z_4\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__22547\,
            I => \sb_translator_1.cntZ0Z_4\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__22544\,
            I => \sb_translator_1.cntZ0Z_4\
        );

    \I__4982\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__22528\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_4\
        );

    \I__4978\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22518\
        );

    \I__4976\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22515\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__22518\,
            I => \N__22512\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__22515\,
            I => mosi_data_out_14
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__22512\,
            I => mosi_data_out_14
        );

    \I__4972\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22503\
        );

    \I__4971\ : InMux
    port map (
            O => \N__22506\,
            I => \N__22499\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22496\
        );

    \I__4969\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22493\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22490\
        );

    \I__4967\ : Odrv12
    port map (
            O => \N__22496\,
            I => \sb_translator_1.cntZ0Z_6\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__22493\,
            I => \sb_translator_1.cntZ0Z_6\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__22490\,
            I => \sb_translator_1.cntZ0Z_6\
        );

    \I__4964\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22477\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__22477\,
            I => \N__22474\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__22474\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_6\
        );

    \I__4960\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__22468\,
            I => \sb_translator_1.state56_a_5_6\
        );

    \I__4958\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__22462\,
            I => \sb_translator_1.state56_a_5_11\
        );

    \I__4956\ : CascadeMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__4955\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__22453\,
            I => \sb_translator_1.state56_a_5_5\
        );

    \I__4953\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__22447\,
            I => \sb_translator_1.state56_a_5_13\
        );

    \I__4951\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22441\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__22441\,
            I => \sb_translator_1.state56_a_5_14\
        );

    \I__4949\ : CascadeMux
    port map (
            O => \N__22438\,
            I => \sb_translator_1.N_318_i_i_o2_12_cascade_\
        );

    \I__4948\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__22429\,
            I => \sb_translator_1.state56_17\
        );

    \I__4945\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22418\
        );

    \I__4943\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22412\
        );

    \I__4942\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22412\
        );

    \I__4941\ : Span4Mux_s3_v
    port map (
            O => \N__22418\,
            I => \N__22409\
        );

    \I__4940\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22406\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__22412\,
            I => \N__22396\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__22409\,
            I => \N__22396\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22393\
        );

    \I__4936\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22382\
        );

    \I__4935\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22382\
        );

    \I__4934\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22382\
        );

    \I__4933\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22382\
        );

    \I__4932\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22382\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__22396\,
            I => \N__22377\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__22393\,
            I => \N__22377\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22374\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__22377\,
            I => \sb_translator_1.state_leds_RNIGMAHZ0\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__22374\,
            I => \sb_translator_1.state_leds_RNIGMAHZ0\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__22369\,
            I => \sb_translator_1.N_318_i_i_o2_15_cascade_\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \sb_translator_1.N_712_cascade_\
        );

    \I__4924\ : CEMux
    port map (
            O => \N__22363\,
            I => \N__22359\
        );

    \I__4923\ : CEMux
    port map (
            O => \N__22362\,
            I => \N__22356\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22350\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22350\
        );

    \I__4920\ : CEMux
    port map (
            O => \N__22355\,
            I => \N__22344\
        );

    \I__4919\ : Span4Mux_v
    port map (
            O => \N__22350\,
            I => \N__22341\
        );

    \I__4918\ : CEMux
    port map (
            O => \N__22349\,
            I => \N__22338\
        );

    \I__4917\ : CEMux
    port map (
            O => \N__22348\,
            I => \N__22327\
        );

    \I__4916\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22315\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22312\
        );

    \I__4914\ : Span4Mux_s0_v
    port map (
            O => \N__22341\,
            I => \N__22307\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__22338\,
            I => \N__22307\
        );

    \I__4912\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22296\
        );

    \I__4911\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22296\
        );

    \I__4910\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22296\
        );

    \I__4909\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22296\
        );

    \I__4908\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22287\
        );

    \I__4907\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22287\
        );

    \I__4906\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22287\
        );

    \I__4905\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22287\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22284\
        );

    \I__4903\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22275\
        );

    \I__4902\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22275\
        );

    \I__4901\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22275\
        );

    \I__4900\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22275\
        );

    \I__4899\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22272\
        );

    \I__4898\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22263\
        );

    \I__4897\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22263\
        );

    \I__4896\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22263\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22263\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__22315\,
            I => \N__22260\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__22312\,
            I => \N__22254\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__22307\,
            I => \N__22254\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22249\
        );

    \I__4890\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22249\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22244\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__22287\,
            I => \N__22244\
        );

    \I__4887\ : Span4Mux_s2_v
    port map (
            O => \N__22284\,
            I => \N__22233\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__22275\,
            I => \N__22233\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22233\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22233\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__22260\,
            I => \N__22233\
        );

    \I__4882\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22230\
        );

    \I__4881\ : Span4Mux_v
    port map (
            O => \N__22254\,
            I => \N__22227\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__22249\,
            I => \N__22220\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__22244\,
            I => \N__22220\
        );

    \I__4878\ : Span4Mux_v
    port map (
            O => \N__22233\,
            I => \N__22220\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22217\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__22227\,
            I => \sb_translator_1.num_leds_1_sqmuxa\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__22220\,
            I => \sb_translator_1.num_leds_1_sqmuxa\
        );

    \I__4874\ : Odrv12
    port map (
            O => \N__22217\,
            I => \sb_translator_1.num_leds_1_sqmuxa\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__22210\,
            I => \N__22207\
        );

    \I__4872\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22193\
        );

    \I__4871\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22176\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22176\
        );

    \I__4869\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22176\
        );

    \I__4868\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22176\
        );

    \I__4867\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22176\
        );

    \I__4866\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22176\
        );

    \I__4865\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22176\
        );

    \I__4864\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22176\
        );

    \I__4863\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22169\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22169\
        );

    \I__4861\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22169\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22166\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__22176\,
            I => \N__22163\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22160\
        );

    \I__4857\ : Span4Mux_v
    port map (
            O => \N__22166\,
            I => \N__22157\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__22163\,
            I => \N__22152\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__22160\,
            I => \N__22152\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__22157\,
            I => \N__22146\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__22152\,
            I => \N__22146\
        );

    \I__4852\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22143\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__22146\,
            I => \N__22140\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__22143\,
            I => \sb_translator_1.stateZ0Z_7\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__22140\,
            I => \sb_translator_1.stateZ0Z_7\
        );

    \I__4848\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__22132\,
            I => \sb_translator_1.state56_a_5_2\
        );

    \I__4846\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__22126\,
            I => \sb_translator_1.state56_a_5_7\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__4843\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__22117\,
            I => \N__22114\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__22114\,
            I => \sb_translator_1.N_318_i_i_o2_0\
        );

    \I__4840\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__22108\,
            I => \sb_translator_1.state56_a_5_12\
        );

    \I__4838\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__22102\,
            I => \sb_translator_1.N_318_i_i_o2_8\
        );

    \I__4836\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__4834\ : Span4Mux_s3_v
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__4832\ : Span4Mux_s3_v
    port map (
            O => \N__22087\,
            I => \N__22084\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__22084\,
            I => \sb_translator_1.N_729\
        );

    \I__4830\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__22078\,
            I => \sb_translator_1.N_712\
        );

    \I__4828\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22067\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__22074\,
            I => \N__22054\
        );

    \I__4826\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22039\
        );

    \I__4825\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22036\
        );

    \I__4824\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22031\
        );

    \I__4823\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22031\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22028\
        );

    \I__4821\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22025\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22018\
        );

    \I__4819\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22018\
        );

    \I__4818\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22018\
        );

    \I__4817\ : InMux
    port map (
            O => \N__22062\,
            I => \N__22010\
        );

    \I__4816\ : InMux
    port map (
            O => \N__22061\,
            I => \N__21998\
        );

    \I__4815\ : InMux
    port map (
            O => \N__22060\,
            I => \N__21998\
        );

    \I__4814\ : InMux
    port map (
            O => \N__22059\,
            I => \N__21998\
        );

    \I__4813\ : InMux
    port map (
            O => \N__22058\,
            I => \N__21998\
        );

    \I__4812\ : InMux
    port map (
            O => \N__22057\,
            I => \N__21998\
        );

    \I__4811\ : InMux
    port map (
            O => \N__22054\,
            I => \N__21984\
        );

    \I__4810\ : InMux
    port map (
            O => \N__22053\,
            I => \N__21984\
        );

    \I__4809\ : InMux
    port map (
            O => \N__22052\,
            I => \N__21977\
        );

    \I__4808\ : InMux
    port map (
            O => \N__22051\,
            I => \N__21977\
        );

    \I__4807\ : InMux
    port map (
            O => \N__22050\,
            I => \N__21977\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22049\,
            I => \N__21966\
        );

    \I__4805\ : InMux
    port map (
            O => \N__22048\,
            I => \N__21966\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22047\,
            I => \N__21966\
        );

    \I__4803\ : InMux
    port map (
            O => \N__22046\,
            I => \N__21966\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22045\,
            I => \N__21966\
        );

    \I__4801\ : InMux
    port map (
            O => \N__22044\,
            I => \N__21959\
        );

    \I__4800\ : InMux
    port map (
            O => \N__22043\,
            I => \N__21959\
        );

    \I__4799\ : InMux
    port map (
            O => \N__22042\,
            I => \N__21959\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__22039\,
            I => \N__21956\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__21945\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__21945\
        );

    \I__4795\ : Span4Mux_v
    port map (
            O => \N__22028\,
            I => \N__21945\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__21945\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__21945\
        );

    \I__4792\ : InMux
    port map (
            O => \N__22017\,
            I => \N__21934\
        );

    \I__4791\ : InMux
    port map (
            O => \N__22016\,
            I => \N__21934\
        );

    \I__4790\ : InMux
    port map (
            O => \N__22015\,
            I => \N__21934\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22014\,
            I => \N__21934\
        );

    \I__4788\ : InMux
    port map (
            O => \N__22013\,
            I => \N__21934\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__21931\
        );

    \I__4786\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21928\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21925\
        );

    \I__4784\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21922\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21905\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21905\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21905\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21905\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21905\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21905\
        );

    \I__4777\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21905\
        );

    \I__4776\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21905\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21898\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21898\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21898\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21891\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__21956\,
            I => \N__21891\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__21945\,
            I => \N__21891\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__21934\,
            I => \N__21884\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__21931\,
            I => \N__21884\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__21928\,
            I => \N__21884\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__21925\,
            I => \N__21881\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21878\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21871\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__21898\,
            I => \N__21871\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__21891\,
            I => \N__21871\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__21884\,
            I => \N__21866\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__21881\,
            I => \N__21866\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__21878\,
            I => \N__21861\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__21871\,
            I => \N__21861\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__21866\,
            I => \sb_translator_1.stateZ0Z_0\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__21861\,
            I => \sb_translator_1.stateZ0Z_0\
        );

    \I__4755\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21852\
        );

    \I__4754\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21849\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21844\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__21849\,
            I => \N__21844\
        );

    \I__4751\ : Span4Mux_v
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__21841\,
            I => \N__21838\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__21838\,
            I => \sb_translator_1.state_RNIOCIR9Z0Z_5\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21832\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21832\,
            I => \sb_translator_1.state56_a_5_4\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21826\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__21826\,
            I => \sb_translator_1.state56_a_5_10\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__4743\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__21817\,
            I => \sb_translator_1.state56_a_5_3\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__21811\,
            I => \sb_translator_1.state56_a_5_16\
        );

    \I__4739\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21805\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__21805\,
            I => \N__21802\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__21799\,
            I => demux_data_in_111
        );

    \I__4735\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__4732\ : Span4Mux_v
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__4731\ : Span4Mux_v
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__21781\,
            I => demux_data_in_39
        );

    \I__4729\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__4727\ : Span4Mux_h
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__4725\ : Odrv4
    port map (
            O => \N__21766\,
            I => demux_data_in_95
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__21763\,
            I => \demux.N_417_i_0_o2Z0Z_0_cascade_\
        );

    \I__4723\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21757\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__21757\,
            I => \demux.N_417_i_0_o2Z0Z_1\
        );

    \I__4721\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21751\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__21751\,
            I => \N__21748\
        );

    \I__4719\ : Span4Mux_v
    port map (
            O => \N__21748\,
            I => \N__21745\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__21745\,
            I => \N__21742\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__21742\,
            I => demux_data_in_47
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__4715\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__21733\,
            I => \demux.N_417_i_0_a3Z0Z_4\
        );

    \I__4713\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__4711\ : Span4Mux_h
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__21721\,
            I => demux_data_in_109
        );

    \I__4709\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__21703\,
            I => demux_data_in_37
        );

    \I__4703\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__21697\,
            I => \N__21694\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__21694\,
            I => \N__21691\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__21691\,
            I => \N__21688\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__21688\,
            I => demux_data_in_93
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__21685\,
            I => \demux.N_419_i_0_o2Z0Z_0_cascade_\
        );

    \I__4697\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__21673\,
            I => \N__21670\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__21670\,
            I => demux_data_in_45
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__21667\,
            I => \demux.N_419_i_0_o2Z0Z_2_cascade_\
        );

    \I__4691\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__21658\,
            I => demux_data_in_13
        );

    \I__4688\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__21652\,
            I => \demux.N_419_i_0_a3Z0Z_5\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__21649\,
            I => \N__21646\
        );

    \I__4685\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__4683\ : Span4Mux_s3_v
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__21634\,
            I => demux_data_in_69
        );

    \I__4680\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__21628\,
            I => \demux.N_419_i_0_a3Z0Z_7\
        );

    \I__4678\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__21622\,
            I => \demux.N_419_i_0_o2Z0Z_8\
        );

    \I__4676\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__21616\,
            I => \N__21611\
        );

    \I__4674\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21608\
        );

    \I__4673\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21605\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__21611\,
            I => \N__21601\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21598\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__21605\,
            I => \N__21595\
        );

    \I__4669\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21592\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__21601\,
            I => \demux.N_422_i_0_o2Z0Z_9\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__21598\,
            I => \demux.N_422_i_0_o2Z0Z_9\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__21595\,
            I => \demux.N_422_i_0_o2Z0Z_9\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__21592\,
            I => \demux.N_422_i_0_o2Z0Z_9\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__21583\,
            I => \N__21580\
        );

    \I__4663\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21571\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__21576\,
            I => \N__21568\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__21575\,
            I => \N__21565\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \N__21562\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__21571\,
            I => \N__21559\
        );

    \I__4657\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21556\
        );

    \I__4656\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21553\
        );

    \I__4655\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21550\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__21559\,
            I => \demux.N_422_i_0_aZ0Z3\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__21556\,
            I => \demux.N_422_i_0_aZ0Z3\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__21553\,
            I => \demux.N_422_i_0_aZ0Z3\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__21550\,
            I => \demux.N_422_i_0_aZ0Z3\
        );

    \I__4650\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__4649\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21532\
        );

    \I__4648\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21529\
        );

    \I__4647\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21526\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__21535\,
            I => \demux.N_422_i_0_o2Z0Z_7\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__21532\,
            I => \demux.N_422_i_0_o2Z0Z_7\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__21529\,
            I => \demux.N_422_i_0_o2Z0Z_7\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__21526\,
            I => \demux.N_422_i_0_o2Z0Z_7\
        );

    \I__4642\ : CEMux
    port map (
            O => \N__21517\,
            I => \N__21513\
        );

    \I__4641\ : CEMux
    port map (
            O => \N__21516\,
            I => \N__21510\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21507\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__21510\,
            I => \N__21504\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__21507\,
            I => \N__21500\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__21504\,
            I => \N__21497\
        );

    \I__4636\ : CEMux
    port map (
            O => \N__21503\,
            I => \N__21494\
        );

    \I__4635\ : Span4Mux_h
    port map (
            O => \N__21500\,
            I => \N__21491\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__21497\,
            I => \N__21488\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21485\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__21491\,
            I => \N__21482\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__21488\,
            I => \N__21479\
        );

    \I__4630\ : Span12Mux_s11_v
    port map (
            O => \N__21485\,
            I => \N__21476\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__21482\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1\
        );

    \I__4628\ : Odrv12
    port map (
            O => \N__21479\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1\
        );

    \I__4627\ : Odrv12
    port map (
            O => \N__21476\,
            I => \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1\
        );

    \I__4626\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21466\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__21466\,
            I => \N__21463\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__21463\,
            I => \N__21460\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__21460\,
            I => mosi_data_out_16
        );

    \I__4622\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21454\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__21454\,
            I => \N__21451\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__21451\,
            I => \N__21448\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__21448\,
            I => \N__21443\
        );

    \I__4618\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21440\
        );

    \I__4617\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21437\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__21443\,
            I => \sb_translator_1.cntZ0Z_8\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__21440\,
            I => \sb_translator_1.cntZ0Z_8\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__21437\,
            I => \sb_translator_1.cntZ0Z_8\
        );

    \I__4613\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21427\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__4611\ : Span4Mux_h
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__21421\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_8\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__21418\,
            I => \N__21413\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__21417\,
            I => \N__21410\
        );

    \I__4607\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21406\
        );

    \I__4606\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21399\
        );

    \I__4605\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21399\
        );

    \I__4604\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21399\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21395\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21392\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21388\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__21395\,
            I => \N__21384\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__21392\,
            I => \N__21381\
        );

    \I__4598\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21378\
        );

    \I__4597\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21373\
        );

    \I__4596\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21373\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__21384\,
            I => \sb_translator_1.cnt_ledsZ0Z_12\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__21381\,
            I => \sb_translator_1.cnt_ledsZ0Z_12\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__21378\,
            I => \sb_translator_1.cnt_ledsZ0Z_12\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__21373\,
            I => \sb_translator_1.cnt_ledsZ0Z_12\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__21364\,
            I => \N__21357\
        );

    \I__4590\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21353\
        );

    \I__4589\ : InMux
    port map (
            O => \N__21362\,
            I => \N__21345\
        );

    \I__4588\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21345\
        );

    \I__4587\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21345\
        );

    \I__4586\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21340\
        );

    \I__4585\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21340\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21337\
        );

    \I__4583\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21334\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__21345\,
            I => \N__21331\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__21340\,
            I => \N__21328\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__21337\,
            I => \N__21325\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__21334\,
            I => \N__21318\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__21331\,
            I => \N__21318\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__21328\,
            I => \N__21318\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__21325\,
            I => \sb_translator_1.cnt_ledsZ0Z_9\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__21318\,
            I => \sb_translator_1.cnt_ledsZ0Z_9\
        );

    \I__4574\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__4573\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21300\
        );

    \I__4572\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21300\
        );

    \I__4571\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21300\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21297\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__21300\,
            I => \N__21294\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__21297\,
            I => \N__21289\
        );

    \I__4567\ : Span4Mux_v
    port map (
            O => \N__21294\,
            I => \N__21289\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__21289\,
            I => \N__21286\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__21286\,
            I => \sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__21283\,
            I => \N__21280\
        );

    \I__4563\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21277\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__21277\,
            I => \N__21274\
        );

    \I__4561\ : Span12Mux_v
    port map (
            O => \N__21274\,
            I => \N__21271\
        );

    \I__4560\ : Odrv12
    port map (
            O => \N__21271\,
            I => demux_data_in_26
        );

    \I__4559\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21265\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__21265\,
            I => \N__21262\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__21262\,
            I => \demux.N_422_i_0_a3Z0Z_7\
        );

    \I__4556\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21256\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__4554\ : Span4Mux_v
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__21250\,
            I => demux_data_in_15
        );

    \I__4552\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21244\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21241\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__21241\,
            I => \N__21238\
        );

    \I__4549\ : Span4Mux_v
    port map (
            O => \N__21238\,
            I => \N__21235\
        );

    \I__4548\ : Span4Mux_v
    port map (
            O => \N__21235\,
            I => \N__21232\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__21232\,
            I => demux_data_in_25
        );

    \I__4546\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21223\
        );

    \I__4544\ : Span4Mux_h
    port map (
            O => \N__21223\,
            I => \N__21220\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__21220\,
            I => demux_data_in_17
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__4541\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21211\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__21211\,
            I => \N__21208\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__21208\,
            I => \N__21205\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__21205\,
            I => demux_data_in_97
        );

    \I__4537\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21196\
        );

    \I__4535\ : Span4Mux_h
    port map (
            O => \N__21196\,
            I => \N__21193\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__4533\ : Odrv4
    port map (
            O => \N__21190\,
            I => demux_data_in_65
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__21187\,
            I => \demux.N_423_i_0_o2Z0Z_4_cascade_\
        );

    \I__4531\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21181\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__21181\,
            I => \demux.N_423_i_0_a3Z0Z_7\
        );

    \I__4529\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21175\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__21175\,
            I => \N__21172\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__21172\,
            I => \N__21169\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__21169\,
            I => \N__21166\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__21166\,
            I => demux_data_in_41
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__21163\,
            I => \demux.N_423_i_0_o2Z0Z_8_cascade_\
        );

    \I__4523\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21157\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__21157\,
            I => \demux.N_423_i_0_o2Z0Z_2\
        );

    \I__4521\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21151\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__21151\,
            I => \demux.N_418_i_0_o2Z0Z_4\
        );

    \I__4519\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21145\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__21145\,
            I => \N__21142\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__21142\,
            I => \N__21139\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__21139\,
            I => \N__21136\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__21136\,
            I => demux_data_in_78
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__21133\,
            I => \demux.N_884_cascade_\
        );

    \I__4513\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21124\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__4510\ : Span4Mux_h
    port map (
            O => \N__21121\,
            I => \N__21118\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__21118\,
            I => demux_data_in_27
        );

    \I__4508\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21112\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__21112\,
            I => \N__21109\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__21109\,
            I => \N__21106\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__21106\,
            I => \N__21103\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__21103\,
            I => demux_data_in_19
        );

    \I__4503\ : CascadeMux
    port map (
            O => \N__21100\,
            I => \N__21097\
        );

    \I__4502\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21094\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21091\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__21091\,
            I => demux_data_in_99
        );

    \I__4499\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21085\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21082\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__21082\,
            I => \N__21079\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__21079\,
            I => \N__21076\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__21076\,
            I => demux_data_in_75
        );

    \I__4494\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21064\
        );

    \I__4493\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21064\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__21071\,
            I => \N__21061\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__21070\,
            I => \N__21056\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__21069\,
            I => \N__21053\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21049\
        );

    \I__4488\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21042\
        );

    \I__4487\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21042\
        );

    \I__4486\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21042\
        );

    \I__4485\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21035\
        );

    \I__4484\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21035\
        );

    \I__4483\ : InMux
    port map (
            O => \N__21052\,
            I => \N__21035\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__21049\,
            I => \N__21030\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__21042\,
            I => \N__21030\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__21035\,
            I => \demux.N_424_i_0_a2Z0Z_0\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__21030\,
            I => \demux.N_424_i_0_a2Z0Z_0\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__21025\,
            I => \demux.N_421_i_0_o2Z0Z_4_cascade_\
        );

    \I__4477\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21019\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__21019\,
            I => \demux.N_421_i_0_a3Z0Z_7\
        );

    \I__4475\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21013\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__21013\,
            I => \N__21010\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__21010\,
            I => \N__21007\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__21007\,
            I => demux_data_in_11
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__21004\,
            I => \demux.N_421_i_0_o2Z0Z_8_cascade_\
        );

    \I__4470\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20998\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__20998\,
            I => \demux.N_421_i_0_o2Z0Z_2\
        );

    \I__4468\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20991\
        );

    \I__4467\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20987\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20984\
        );

    \I__4465\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20981\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20977\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20972\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20972\
        );

    \I__4461\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20969\
        );

    \I__4460\ : Odrv4
    port map (
            O => \N__20977\,
            I => \demux.N_422_i_0_o2Z0Z_8\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__20972\,
            I => \demux.N_422_i_0_o2Z0Z_8\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__20969\,
            I => \demux.N_422_i_0_o2Z0Z_8\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__20962\,
            I => \N__20958\
        );

    \I__4456\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20953\
        );

    \I__4455\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20953\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20950\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__20950\,
            I => \N__20943\
        );

    \I__4452\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20940\
        );

    \I__4451\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20937\
        );

    \I__4450\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20932\
        );

    \I__4449\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20932\
        );

    \I__4448\ : Span4Mux_h
    port map (
            O => \N__20943\,
            I => \N__20929\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__20940\,
            I => \sb_translator_1.num_ledsZ0Z_15\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__20937\,
            I => \sb_translator_1.num_ledsZ0Z_15\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__20932\,
            I => \sb_translator_1.num_ledsZ0Z_15\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__20929\,
            I => \sb_translator_1.num_ledsZ0Z_15\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__20920\,
            I => \N__20917\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20913\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20910\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__20913\,
            I => \sb_translator_1.cnt_leds_i_16\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__20910\,
            I => \sb_translator_1.cnt_leds_i_16\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20900\
        );

    \I__4437\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20895\
        );

    \I__4436\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20895\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__20900\,
            I => \sb_translator_1.cnt_ledsZ0Z_15\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__20895\,
            I => \sb_translator_1.cnt_ledsZ0Z_15\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__4432\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20884\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20881\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__20881\,
            I => \sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15\
        );

    \I__4429\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20871\
        );

    \I__4428\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20871\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__20876\,
            I => \N__20867\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20862\
        );

    \I__4425\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20857\
        );

    \I__4424\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20857\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20852\
        );

    \I__4422\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20852\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__20862\,
            I => \N__20849\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__20857\,
            I => \sb_translator_1.num_ledsZ0Z_12\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__20852\,
            I => \sb_translator_1.num_ledsZ0Z_12\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__20849\,
            I => \sb_translator_1.num_ledsZ0Z_12\
        );

    \I__4417\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20837\
        );

    \I__4416\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20832\
        );

    \I__4415\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20832\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__20837\,
            I => \sb_translator_1.cnt_ledsZ0Z_13\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__20832\,
            I => \sb_translator_1.cnt_ledsZ0Z_13\
        );

    \I__4412\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20824\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__4410\ : Span4Mux_s3_v
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__20818\,
            I => \sb_translator_1.cnt_leds_RNI15HTZ0Z_13\
        );

    \I__4408\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20803\
        );

    \I__4407\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20803\
        );

    \I__4406\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20803\
        );

    \I__4405\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20803\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20799\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20795\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__20799\,
            I => \N__20792\
        );

    \I__4401\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20787\
        );

    \I__4400\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20787\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__20792\,
            I => \sb_translator_1.num_ledsZ0Z_14\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__20787\,
            I => \sb_translator_1.num_ledsZ0Z_14\
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__20782\,
            I => \N__20777\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20766\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20766\
        );

    \I__4394\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20766\
        );

    \I__4393\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20766\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__20775\,
            I => \N__20762\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__20766\,
            I => \N__20759\
        );

    \I__4390\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20754\
        );

    \I__4389\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20754\
        );

    \I__4388\ : Span4Mux_h
    port map (
            O => \N__20759\,
            I => \N__20751\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__20754\,
            I => \sb_translator_1.num_ledsZ0Z_13\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__20751\,
            I => \sb_translator_1.num_ledsZ0Z_13\
        );

    \I__4385\ : CascadeMux
    port map (
            O => \N__20746\,
            I => \sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_\
        );

    \I__4384\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20738\
        );

    \I__4383\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20733\
        );

    \I__4382\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20733\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__20738\,
            I => \sb_translator_1.cnt_ledsZ0Z_14\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__20733\,
            I => \sb_translator_1.cnt_ledsZ0Z_14\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__20728\,
            I => \N__20725\
        );

    \I__4378\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__20719\,
            I => \sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__4374\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__4372\ : Span12Mux_s11_v
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__4371\ : Odrv12
    port map (
            O => \N__20704\,
            I => demux_data_in_66
        );

    \I__4370\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20695\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__20695\,
            I => \N__20692\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__20692\,
            I => \N__20689\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__20689\,
            I => demux_data_in_30
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__20686\,
            I => \N__20683\
        );

    \I__4364\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20677\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__20677\,
            I => demux_data_in_102
        );

    \I__4361\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__20671\,
            I => \N__20668\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__20665\,
            I => \N__20662\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__20662\,
            I => demux_data_in_32
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__4355\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__20650\,
            I => \N__20647\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__20647\,
            I => demux_data_in_104
        );

    \I__4351\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__20641\,
            I => \demux.N_424_i_0_o2_0Z0Z_0\
        );

    \I__4349\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__20632\,
            I => \N__20629\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__20626\,
            I => demux_data_in_44
        );

    \I__4344\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20620\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__20620\,
            I => \N__20617\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__20617\,
            I => \N__20614\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__20614\,
            I => \N__20611\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__20611\,
            I => demux_data_in_22
        );

    \I__4339\ : InMux
    port map (
            O => \N__20608\,
            I => \sb_translator_1.state56_a_5_cry_12\
        );

    \I__4338\ : InMux
    port map (
            O => \N__20605\,
            I => \sb_translator_1.state56_a_5_cry_13\
        );

    \I__4337\ : InMux
    port map (
            O => \N__20602\,
            I => \bfn_8_5_0_\
        );

    \I__4336\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20595\
        );

    \I__4335\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20592\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__20595\,
            I => \sb_translator_1.cnt_ledsZ0Z_16\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__20592\,
            I => \sb_translator_1.cnt_ledsZ0Z_16\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__20587\,
            I => \sb_translator_1.cnt_leds_i_16_cascade_\
        );

    \I__4331\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__20578\,
            I => \sb_translator_1.num_leds_RNIOJBMZ0Z_15\
        );

    \I__4328\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20571\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__20574\,
            I => \N__20568\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__20571\,
            I => \N__20565\
        );

    \I__4325\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20562\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__20565\,
            I => \N__20557\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20557\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__20557\,
            I => \sb_translator_1.num_leds_RNIU1HTZ0Z_11\
        );

    \I__4321\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20551\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20548\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__20548\,
            I => \sb_translator_1.cnt_leds_RNIV62R1Z0Z_13\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__20545\,
            I => \N__20542\
        );

    \I__4317\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20539\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20536\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__20536\,
            I => \sb_translator_1.cnt_leds_RNI48HTZ0Z_14\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__20533\,
            I => \sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_\
        );

    \I__4313\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20527\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20524\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__20524\,
            I => \sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15\
        );

    \I__4310\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__20518\,
            I => \sb_translator_1.cnt_leds_RNIHCUTZ0Z_7\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__20515\,
            I => \N__20512\
        );

    \I__4307\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__20509\,
            I => \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6\
        );

    \I__4305\ : InMux
    port map (
            O => \N__20506\,
            I => \sb_translator_1.state56_a_5_cry_4\
        );

    \I__4304\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__20500\,
            I => \sb_translator_1.cnt_leds_RNINIUTZ0Z_8\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__20497\,
            I => \N__20494\
        );

    \I__4301\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__20491\,
            I => \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7\
        );

    \I__4299\ : InMux
    port map (
            O => \N__20488\,
            I => \sb_translator_1.state56_a_5_cry_5\
        );

    \I__4298\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__20479\,
            I => \sb_translator_1.num_leds_RNITOUTZ0Z_8\
        );

    \I__4295\ : InMux
    port map (
            O => \N__20476\,
            I => \N__20472\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__20475\,
            I => \N__20469\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20466\
        );

    \I__4292\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20463\
        );

    \I__4291\ : Span4Mux_v
    port map (
            O => \N__20466\,
            I => \N__20460\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20457\
        );

    \I__4289\ : Odrv4
    port map (
            O => \N__20460\,
            I => \sb_translator_1.cnt_leds_RNITAVEZ0Z_8\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__20457\,
            I => \sb_translator_1.cnt_leds_RNITAVEZ0Z_8\
        );

    \I__4287\ : InMux
    port map (
            O => \N__20452\,
            I => \bfn_8_4_0_\
        );

    \I__4286\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__20443\,
            I => \sb_translator_1.num_leds_RNIH2E91Z0Z_9\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__4282\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20433\
        );

    \I__4281\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20430\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20427\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__20430\,
            I => \sb_translator_1.num_leds_RNI0EVEZ0Z_8\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__20427\,
            I => \sb_translator_1.num_leds_RNI0EVEZ0Z_8\
        );

    \I__4277\ : InMux
    port map (
            O => \N__20422\,
            I => \sb_translator_1.state56_a_5_cry_7\
        );

    \I__4276\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__20413\,
            I => \sb_translator_1.num_leds_RNICJVN1Z0Z_10\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__20410\,
            I => \N__20407\
        );

    \I__4272\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__20404\,
            I => \N__20401\
        );

    \I__4270\ : Odrv12
    port map (
            O => \N__20401\,
            I => \sb_translator_1.num_leds_RNIHKEQZ0Z_9\
        );

    \I__4269\ : InMux
    port map (
            O => \N__20398\,
            I => \sb_translator_1.state56_a_5_cry_8\
        );

    \I__4268\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__20389\,
            I => \sb_translator_1.num_leds_RNIP02R1Z0Z_11\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__4264\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__20380\,
            I => \N__20377\
        );

    \I__4262\ : Odrv12
    port map (
            O => \N__20377\,
            I => \sb_translator_1.num_leds_RNIRUGTZ0Z_10\
        );

    \I__4261\ : InMux
    port map (
            O => \N__20374\,
            I => \sb_translator_1.state56_a_5_cry_9\
        );

    \I__4260\ : InMux
    port map (
            O => \N__20371\,
            I => \sb_translator_1.state56_a_5_cry_10\
        );

    \I__4259\ : InMux
    port map (
            O => \N__20368\,
            I => \sb_translator_1.state56_a_5_cry_11\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__4257\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20355\
        );

    \I__4256\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20348\
        );

    \I__4255\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20348\
        );

    \I__4254\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20348\
        );

    \I__4253\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20345\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20342\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__20348\,
            I => \N__20339\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20336\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__20342\,
            I => \N__20333\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__20339\,
            I => \N__20330\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__20336\,
            I => \N__20327\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__20333\,
            I => ram_sel_13
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__20330\,
            I => ram_sel_13
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__20327\,
            I => ram_sel_13
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__20320\,
            I => \N__20313\
        );

    \I__4242\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20309\
        );

    \I__4241\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20302\
        );

    \I__4240\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20302\
        );

    \I__4239\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20302\
        );

    \I__4238\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20297\
        );

    \I__4237\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20297\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__20309\,
            I => \N__20294\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20291\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20288\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__20294\,
            I => \N__20283\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__20291\,
            I => \N__20283\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__20288\,
            I => \N__20280\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__20283\,
            I => ram_sel_10
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__20280\,
            I => ram_sel_10
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \N__20270\
        );

    \I__4227\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20264\
        );

    \I__4226\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20259\
        );

    \I__4225\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20259\
        );

    \I__4224\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20254\
        );

    \I__4223\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20254\
        );

    \I__4222\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20251\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__20264\,
            I => \N__20246\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__20259\,
            I => \N__20246\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__20254\,
            I => \N__20243\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20240\
        );

    \I__4217\ : Span4Mux_h
    port map (
            O => \N__20246\,
            I => \N__20237\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__20243\,
            I => \N__20234\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__20240\,
            I => ram_sel_7
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__20237\,
            I => ram_sel_7
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__20234\,
            I => ram_sel_7
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__20227\,
            I => \N__20223\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__20226\,
            I => \N__20218\
        );

    \I__4210\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20212\
        );

    \I__4209\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20212\
        );

    \I__4208\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20209\
        );

    \I__4207\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20204\
        );

    \I__4206\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20204\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__20212\,
            I => \demux.N_240\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__20209\,
            I => \demux.N_240\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20204\,
            I => \demux.N_240\
        );

    \I__4202\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20194\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__20194\,
            I => \N__20191\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__20185\,
            I => \N__20182\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__20182\,
            I => demux_data_in_29
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__20179\,
            I => \N__20176\
        );

    \I__4195\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20173\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__20173\,
            I => \N__20169\
        );

    \I__4193\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20166\
        );

    \I__4192\ : Span4Mux_s2_v
    port map (
            O => \N__20169\,
            I => \N__20161\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__20166\,
            I => \N__20161\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__20161\,
            I => \sb_translator_1.state56_a_5_ac0_1\
        );

    \I__4189\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__20155\,
            I => \sb_translator_1.cnt_leds_RNIJDTTZ0Z_2\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__20152\,
            I => \N__20149\
        );

    \I__4186\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__20146\,
            I => \sb_translator_1.state56_a_5_44\
        );

    \I__4184\ : InMux
    port map (
            O => \N__20143\,
            I => \sb_translator_1.state56_a_5_cry_0_c_THRU_CO\
        );

    \I__4183\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20137\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__20137\,
            I => \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__20134\,
            I => \N__20131\
        );

    \I__4180\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20128\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__20128\,
            I => \sb_translator_1.cnt_leds_RNIPJTTZ0Z_3\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20125\,
            I => \sb_translator_1.state56_a_5_cry_0\
        );

    \I__4177\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__20119\,
            I => \sb_translator_1.cnt_leds_RNIERUEZ0Z_3\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20113\
        );

    \I__4174\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__20110\,
            I => \sb_translator_1.cnt_leds_RNIVPTTZ0Z_4\
        );

    \I__4172\ : InMux
    port map (
            O => \N__20107\,
            I => \sb_translator_1.state56_a_5_cry_1\
        );

    \I__4171\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20100\
        );

    \I__4170\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20097\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__20100\,
            I => \sb_translator_1.cnt_leds_RNIHUUEZ0Z_4\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__20097\,
            I => \sb_translator_1.cnt_leds_RNIHUUEZ0Z_4\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__4166\ : InMux
    port map (
            O => \N__20089\,
            I => \N__20086\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__20086\,
            I => \sb_translator_1.cnt_leds_RNI50UTZ0Z_5\
        );

    \I__4164\ : InMux
    port map (
            O => \N__20083\,
            I => \sb_translator_1.state56_a_5_cry_2\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20077\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__20077\,
            I => \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__20074\,
            I => \N__20071\
        );

    \I__4160\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20068\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__20068\,
            I => \sb_translator_1.cnt_leds_RNIB6UTZ0Z_6\
        );

    \I__4158\ : InMux
    port map (
            O => \N__20065\,
            I => \sb_translator_1.state56_a_5_cry_3\
        );

    \I__4157\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20059\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__20059\,
            I => \demux.N_917\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__20056\,
            I => \demux.N_424_i_0_o2_0_7_cascade_\
        );

    \I__4154\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__20050\,
            I => \demux.N_424_i_0_o2_0_10\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__20047\,
            I => \demux.N_424_i_0_o2Z0Z_0_cascade_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20041\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__20041\,
            I => \N__20038\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__20038\,
            I => \N__20035\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__20035\,
            I => demux_data_in_16
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__20032\,
            I => \N__20029\
        );

    \I__4146\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__20023\,
            I => \N__20020\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__20020\,
            I => demux_data_in_96
        );

    \I__4142\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__20011\,
            I => \N__20008\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__20008\,
            I => demux_data_in_64
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__20005\,
            I => \demux.N_424_i_0_o2Z0Z_4_cascade_\
        );

    \I__4137\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19998\
        );

    \I__4136\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19995\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19991\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__19995\,
            I => \N__19988\
        );

    \I__4133\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19985\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__19991\,
            I => \N__19978\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__19988\,
            I => \N__19978\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19978\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__19978\,
            I => \demux.N_424_i_0_o2Z0Z_8\
        );

    \I__4128\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19967\
        );

    \I__4126\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19964\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__19970\,
            I => \N__19961\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__19967\,
            I => \N__19956\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19956\
        );

    \I__4122\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19953\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__19956\,
            I => \demux.N_424_i_0_aZ0Z3\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__19953\,
            I => \demux.N_424_i_0_aZ0Z3\
        );

    \I__4119\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19944\
        );

    \I__4118\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19941\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__19944\,
            I => \N__19937\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19934\
        );

    \I__4115\ : InMux
    port map (
            O => \N__19940\,
            I => \N__19931\
        );

    \I__4114\ : Span4Mux_h
    port map (
            O => \N__19937\,
            I => \N__19925\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__19934\,
            I => \N__19925\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19922\
        );

    \I__4111\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19919\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__19925\,
            I => \demux.N_424_i_0_o2_9\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__19922\,
            I => \demux.N_424_i_0_o2_9\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__19919\,
            I => \demux.N_424_i_0_o2_9\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__19912\,
            I => \demux.N_424_i_0_o2Z0Z_8_cascade_\
        );

    \I__4106\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19905\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__19908\,
            I => \N__19902\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__19905\,
            I => \N__19899\
        );

    \I__4103\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19896\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__19899\,
            I => \N__19889\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19889\
        );

    \I__4100\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19886\
        );

    \I__4099\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19883\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__19889\,
            I => \demux.N_424_i_0_o2Z0Z_7\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__19886\,
            I => \demux.N_424_i_0_o2Z0Z_7\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__19883\,
            I => \demux.N_424_i_0_o2Z0Z_7\
        );

    \I__4095\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19873\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19870\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__4091\ : Span4Mux_v
    port map (
            O => \N__19864\,
            I => \N__19861\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__19861\,
            I => demux_data_in_24
        );

    \I__4089\ : InMux
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__19855\,
            I => \demux.N_424_i_0_a3Z0Z_7\
        );

    \I__4087\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19849\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__19849\,
            I => \N__19845\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__19848\,
            I => \N__19841\
        );

    \I__4084\ : Span4Mux_v
    port map (
            O => \N__19845\,
            I => \N__19837\
        );

    \I__4083\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19834\
        );

    \I__4082\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19831\
        );

    \I__4081\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19828\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__19837\,
            I => ram_sel_0
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__19834\,
            I => ram_sel_0
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__19831\,
            I => ram_sel_0
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__19828\,
            I => ram_sel_0
        );

    \I__4076\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19814\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \N__19811\
        );

    \I__4074\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19807\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__19814\,
            I => \N__19803\
        );

    \I__4072\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19798\
        );

    \I__4071\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19798\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19795\
        );

    \I__4069\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19792\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__19803\,
            I => \N__19789\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19786\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__19795\,
            I => \N__19783\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__19792\,
            I => \N__19780\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__19789\,
            I => ram_sel_11
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__19786\,
            I => ram_sel_11
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__19783\,
            I => ram_sel_11
        );

    \I__4061\ : Odrv12
    port map (
            O => \N__19780\,
            I => ram_sel_11
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__19771\,
            I => \demux.N_906_cascade_\
        );

    \I__4059\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19764\
        );

    \I__4058\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19761\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__19764\,
            I => \N__19758\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19753\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__19758\,
            I => \N__19749\
        );

    \I__4054\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19744\
        );

    \I__4053\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19744\
        );

    \I__4052\ : Span4Mux_h
    port map (
            O => \N__19753\,
            I => \N__19741\
        );

    \I__4051\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19738\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__19749\,
            I => ram_sel_4
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__19744\,
            I => ram_sel_4
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__19741\,
            I => ram_sel_4
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__19738\,
            I => ram_sel_4
        );

    \I__4046\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19726\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__19726\,
            I => \demux.N_424_i_0_o2_0Z0Z_3\
        );

    \I__4044\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19717\
        );

    \I__4042\ : Span4Mux_v
    port map (
            O => \N__19717\,
            I => \N__19714\
        );

    \I__4041\ : Span4Mux_h
    port map (
            O => \N__19714\,
            I => \N__19711\
        );

    \I__4040\ : Span4Mux_v
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__19708\,
            I => demux_data_in_28
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__19705\,
            I => \demux.N_918_cascade_\
        );

    \I__4037\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19699\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__19699\,
            I => \N__19696\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__19693\,
            I => demux_data_in_105
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__19690\,
            I => \demux.N_424_i_0_a2Z0Z_5_cascade_\
        );

    \I__4032\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__19675\,
            I => demux_data_in_33
        );

    \I__4027\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19669\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__19669\,
            I => \demux.N_423_i_0_o2Z0Z_0\
        );

    \I__4025\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19662\
        );

    \I__4024\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19659\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__19662\,
            I => \demux.N_918\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__19659\,
            I => \demux.N_918\
        );

    \I__4021\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19646\
        );

    \I__4020\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19646\
        );

    \I__4019\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19637\
        );

    \I__4018\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19637\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19634\
        );

    \I__4016\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19625\
        );

    \I__4015\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19625\
        );

    \I__4014\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19625\
        );

    \I__4013\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19625\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__19637\,
            I => \N__19618\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__19634\,
            I => \N__19618\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19618\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__19618\,
            I => \demux.N_424_i_0_a2Z0Z_7\
        );

    \I__4008\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19612\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__19612\,
            I => \N__19609\
        );

    \I__4006\ : Span4Mux_h
    port map (
            O => \N__19609\,
            I => \N__19606\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__19606\,
            I => \demux.N_424_i_0_o2_0_1\
        );

    \I__4004\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19599\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__19602\,
            I => \N__19596\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__19599\,
            I => \N__19592\
        );

    \I__4001\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19587\
        );

    \I__4000\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19587\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__19592\,
            I => \N__19584\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19579\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__19584\,
            I => \N__19579\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__19579\,
            I => \demux.N_236\
        );

    \I__3995\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19573\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__19573\,
            I => \N__19570\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__19570\,
            I => \N__19566\
        );

    \I__3992\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19563\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__19566\,
            I => \demux.N_235\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__19563\,
            I => \demux.N_235\
        );

    \I__3989\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19555\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__19555\,
            I => \demux.N_424_i_0_o2_0Z0Z_2\
        );

    \I__3987\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19547\
        );

    \I__3986\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19542\
        );

    \I__3985\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19542\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__19547\,
            I => \demux.N_237\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__19542\,
            I => \demux.N_237\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__19537\,
            I => \demux.N_424_i_0_o2_0_8Z0Z_1_cascade_\
        );

    \I__3981\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19529\
        );

    \I__3980\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19524\
        );

    \I__3979\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19524\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__19529\,
            I => \demux.N_238\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__19524\,
            I => \demux.N_238\
        );

    \I__3976\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__19510\,
            I => demux_data_in_91
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__19507\,
            I => \demux.N_421_i_0_o2Z0Z_0_cascade_\
        );

    \I__3971\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__19498\,
            I => \N__19495\
        );

    \I__3968\ : Span4Mux_h
    port map (
            O => \N__19495\,
            I => \N__19492\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__19492\,
            I => demux_data_in_2
        );

    \I__3966\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__3964\ : Span4Mux_v
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__19480\,
            I => demux_data_in_106
        );

    \I__3962\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__19468\,
            I => demux_data_in_34
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__19465\,
            I => \demux.N_422_i_0_o2Z0Z_0_cascade_\
        );

    \I__3957\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19459\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__3955\ : Span4Mux_v
    port map (
            O => \N__19456\,
            I => \N__19453\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__19453\,
            I => demux_data_in_90
        );

    \I__3953\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19447\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__19447\,
            I => \demux.N_422_i_0_a3Z0Z_4\
        );

    \I__3951\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19441\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__19435\,
            I => demux_data_in_10
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \demux.N_422_i_0_o2Z0Z_1_cascade_\
        );

    \I__3946\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19423\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__19420\,
            I => demux_data_in_9
        );

    \I__3942\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19414\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__19411\,
            I => \N__19408\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__19408\,
            I => demux_data_in_89
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__19405\,
            I => \demux.N_423_i_0_a3Z0Z_5_cascade_\
        );

    \I__3937\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__19393\,
            I => demux_data_in_43
        );

    \I__3933\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__19387\,
            I => \demux.N_837\
        );

    \I__3931\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19380\
        );

    \I__3930\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19377\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__19380\,
            I => \demux.N_424_i_0_a2Z0Z_34\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__19377\,
            I => \demux.N_424_i_0_a2Z0Z_34\
        );

    \I__3927\ : InMux
    port map (
            O => \N__19372\,
            I => \sb_translator_1.cnt_leds_cry_14\
        );

    \I__3926\ : InMux
    port map (
            O => \N__19369\,
            I => \bfn_7_6_0_\
        );

    \I__3925\ : CEMux
    port map (
            O => \N__19366\,
            I => \N__19362\
        );

    \I__3924\ : CEMux
    port map (
            O => \N__19365\,
            I => \N__19359\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__19362\,
            I => \N__19356\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19352\
        );

    \I__3921\ : Span4Mux_v
    port map (
            O => \N__19356\,
            I => \N__19349\
        );

    \I__3920\ : CEMux
    port map (
            O => \N__19355\,
            I => \N__19346\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__19352\,
            I => \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__19349\,
            I => \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__19346\,
            I => \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1\
        );

    \I__3916\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19336\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19333\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__19333\,
            I => \N__19330\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__19330\,
            I => demux_data_in_40
        );

    \I__3912\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__3910\ : Span4Mux_v
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__19318\,
            I => demux_data_in_88
        );

    \I__3908\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19312\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__19312\,
            I => \demux.N_424_i_0_a3Z0Z_4\
        );

    \I__3906\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19303\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__19303\,
            I => \N__19300\
        );

    \I__3903\ : Span4Mux_v
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__19297\,
            I => demux_data_in_8
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__19294\,
            I => \demux.N_424_i_0_o2Z0Z_1_cascade_\
        );

    \I__3900\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19285\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__19285\,
            I => \N__19282\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__19282\,
            I => \N__19279\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__19279\,
            I => demux_data_in_0
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__19276\,
            I => \demux.N_424_i_0_aZ0Z3_cascade_\
        );

    \I__3894\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19270\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__19264\,
            I => demux_data_in_35
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__3889\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19255\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19252\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__19252\,
            I => \N__19249\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__19249\,
            I => demux_data_in_107
        );

    \I__3885\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19238\
        );

    \I__3884\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19238\
        );

    \I__3883\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19235\
        );

    \I__3882\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19232\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19229\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__19235\,
            I => \sb_translator_1.cnt_ledsZ0Z_7\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__19232\,
            I => \sb_translator_1.cnt_ledsZ0Z_7\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__19229\,
            I => \sb_translator_1.cnt_ledsZ0Z_7\
        );

    \I__3877\ : InMux
    port map (
            O => \N__19222\,
            I => \sb_translator_1.cnt_leds_cry_6\
        );

    \I__3876\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19216\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__19216\,
            I => \N__19210\
        );

    \I__3874\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19205\
        );

    \I__3873\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19205\
        );

    \I__3872\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19202\
        );

    \I__3871\ : Sp12to4
    port map (
            O => \N__19210\,
            I => \N__19197\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19197\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__19202\,
            I => \sb_translator_1.cnt_ledsZ0Z_8\
        );

    \I__3868\ : Odrv12
    port map (
            O => \N__19197\,
            I => \sb_translator_1.cnt_ledsZ0Z_8\
        );

    \I__3867\ : InMux
    port map (
            O => \N__19192\,
            I => \bfn_7_5_0_\
        );

    \I__3866\ : InMux
    port map (
            O => \N__19189\,
            I => \sb_translator_1.cnt_leds_cry_8\
        );

    \I__3865\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19177\
        );

    \I__3864\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19172\
        );

    \I__3863\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19172\
        );

    \I__3862\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19163\
        );

    \I__3861\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19163\
        );

    \I__3860\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19163\
        );

    \I__3859\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19163\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__19177\,
            I => \sb_translator_1.cnt_ledsZ0Z_10\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__19172\,
            I => \sb_translator_1.cnt_ledsZ0Z_10\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__19163\,
            I => \sb_translator_1.cnt_ledsZ0Z_10\
        );

    \I__3855\ : InMux
    port map (
            O => \N__19156\,
            I => \sb_translator_1.cnt_leds_cry_9\
        );

    \I__3854\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19144\
        );

    \I__3853\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19141\
        );

    \I__3852\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19138\
        );

    \I__3851\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19129\
        );

    \I__3850\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19129\
        );

    \I__3849\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19129\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19129\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__19144\,
            I => \sb_translator_1.cnt_ledsZ0Z_11\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__19141\,
            I => \sb_translator_1.cnt_ledsZ0Z_11\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__19138\,
            I => \sb_translator_1.cnt_ledsZ0Z_11\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__19129\,
            I => \sb_translator_1.cnt_ledsZ0Z_11\
        );

    \I__3843\ : InMux
    port map (
            O => \N__19120\,
            I => \sb_translator_1.cnt_leds_cry_10\
        );

    \I__3842\ : InMux
    port map (
            O => \N__19117\,
            I => \sb_translator_1.cnt_leds_cry_11\
        );

    \I__3841\ : InMux
    port map (
            O => \N__19114\,
            I => \sb_translator_1.cnt_leds_cry_12\
        );

    \I__3840\ : InMux
    port map (
            O => \N__19111\,
            I => \sb_translator_1.cnt_leds_cry_13\
        );

    \I__3839\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19101\
        );

    \I__3837\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19098\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__19101\,
            I => \N__19090\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19090\
        );

    \I__3834\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19085\
        );

    \I__3833\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19085\
        );

    \I__3832\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19082\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__19090\,
            I => \sb_translator_1.cnt19\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__19085\,
            I => \sb_translator_1.cnt19\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__19082\,
            I => \sb_translator_1.cnt19\
        );

    \I__3828\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19062\
        );

    \I__3827\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19062\
        );

    \I__3826\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19062\
        );

    \I__3825\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19062\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__19071\,
            I => \N__19058\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19055\
        );

    \I__3822\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19050\
        );

    \I__3821\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19050\
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__19055\,
            I => \sb_translator_1.num_ledsZ0Z_2\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__19050\,
            I => \sb_translator_1.num_ledsZ0Z_2\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \sb_translator_1.state56_a_5_44_cascade_\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \N__19038\
        );

    \I__3816\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19030\
        );

    \I__3815\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19030\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__19037\,
            I => \N__19027\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19024\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__19035\,
            I => \N__19020\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__19030\,
            I => \N__19016\
        );

    \I__3810\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19013\
        );

    \I__3809\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19004\
        );

    \I__3808\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19004\
        );

    \I__3807\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19004\
        );

    \I__3806\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19004\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__19016\,
            I => \sb_translator_1.num_ledsZ0Z_1\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__19013\,
            I => \sb_translator_1.num_ledsZ0Z_1\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__19004\,
            I => \sb_translator_1.num_ledsZ0Z_1\
        );

    \I__3802\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__3801\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18988\
        );

    \I__3800\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18985\
        );

    \I__3799\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18982\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__18991\,
            I => \sb_translator_1.cnt_ledsZ0Z_0\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18988\,
            I => \sb_translator_1.cnt_ledsZ0Z_0\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__18985\,
            I => \sb_translator_1.cnt_ledsZ0Z_0\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__18982\,
            I => \sb_translator_1.cnt_ledsZ0Z_0\
        );

    \I__3794\ : InMux
    port map (
            O => \N__18973\,
            I => \bfn_7_4_0_\
        );

    \I__3793\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18963\
        );

    \I__3792\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18960\
        );

    \I__3791\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18955\
        );

    \I__3790\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18955\
        );

    \I__3789\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18952\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__18963\,
            I => \sb_translator_1.cnt_ledsZ0Z_1\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__18960\,
            I => \sb_translator_1.cnt_ledsZ0Z_1\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18955\,
            I => \sb_translator_1.cnt_ledsZ0Z_1\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__18952\,
            I => \sb_translator_1.cnt_ledsZ0Z_1\
        );

    \I__3784\ : InMux
    port map (
            O => \N__18943\,
            I => \sb_translator_1.cnt_leds_cry_0\
        );

    \I__3783\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18931\
        );

    \I__3781\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18926\
        );

    \I__3780\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18926\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__18934\,
            I => \sb_translator_1.cnt_ledsZ0Z_2\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__18931\,
            I => \sb_translator_1.cnt_ledsZ0Z_2\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__18926\,
            I => \sb_translator_1.cnt_ledsZ0Z_2\
        );

    \I__3776\ : InMux
    port map (
            O => \N__18919\,
            I => \sb_translator_1.cnt_leds_cry_1\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__18916\,
            I => \N__18911\
        );

    \I__3774\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18907\
        );

    \I__3773\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18904\
        );

    \I__3772\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18899\
        );

    \I__3771\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18899\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__18907\,
            I => \sb_translator_1.cnt_ledsZ0Z_3\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__18904\,
            I => \sb_translator_1.cnt_ledsZ0Z_3\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__18899\,
            I => \sb_translator_1.cnt_ledsZ0Z_3\
        );

    \I__3767\ : InMux
    port map (
            O => \N__18892\,
            I => \sb_translator_1.cnt_leds_cry_2\
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__18889\,
            I => \N__18884\
        );

    \I__3765\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18880\
        );

    \I__3764\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18877\
        );

    \I__3763\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18872\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18872\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__18880\,
            I => \sb_translator_1.cnt_ledsZ0Z_4\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__18877\,
            I => \sb_translator_1.cnt_ledsZ0Z_4\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__18872\,
            I => \sb_translator_1.cnt_ledsZ0Z_4\
        );

    \I__3758\ : InMux
    port map (
            O => \N__18865\,
            I => \sb_translator_1.cnt_leds_cry_3\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__18862\,
            I => \N__18859\
        );

    \I__3756\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18851\
        );

    \I__3755\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18851\
        );

    \I__3754\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18848\
        );

    \I__3753\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18845\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__18851\,
            I => \N__18842\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__18848\,
            I => \sb_translator_1.cnt_ledsZ0Z_5\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__18845\,
            I => \sb_translator_1.cnt_ledsZ0Z_5\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__18842\,
            I => \sb_translator_1.cnt_ledsZ0Z_5\
        );

    \I__3748\ : InMux
    port map (
            O => \N__18835\,
            I => \sb_translator_1.cnt_leds_cry_4\
        );

    \I__3747\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18824\
        );

    \I__3746\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18824\
        );

    \I__3745\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18821\
        );

    \I__3744\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18818\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__18824\,
            I => \N__18815\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__18821\,
            I => \sb_translator_1.cnt_ledsZ0Z_6\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__18818\,
            I => \sb_translator_1.cnt_ledsZ0Z_6\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__18815\,
            I => \sb_translator_1.cnt_ledsZ0Z_6\
        );

    \I__3739\ : InMux
    port map (
            O => \N__18808\,
            I => \sb_translator_1.cnt_leds_cry_5\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__18805\,
            I => \N__18801\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__18804\,
            I => \N__18797\
        );

    \I__3736\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18786\
        );

    \I__3735\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18786\
        );

    \I__3734\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18786\
        );

    \I__3733\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18786\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__18795\,
            I => \N__18782\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__18786\,
            I => \N__18779\
        );

    \I__3730\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18774\
        );

    \I__3729\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18774\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__18779\,
            I => \sb_translator_1.num_ledsZ0Z_6\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__18774\,
            I => \sb_translator_1.num_ledsZ0Z_6\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__18769\,
            I => \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_\
        );

    \I__3725\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18754\
        );

    \I__3724\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18754\
        );

    \I__3723\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18754\
        );

    \I__3722\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18754\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18750\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__18753\,
            I => \N__18746\
        );

    \I__3719\ : Span4Mux_s2_v
    port map (
            O => \N__18750\,
            I => \N__18743\
        );

    \I__3718\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18738\
        );

    \I__3717\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18738\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__18743\,
            I => \sb_translator_1.num_ledsZ0Z_7\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__18738\,
            I => \sb_translator_1.num_ledsZ0Z_7\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18730\
        );

    \I__3713\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18723\
        );

    \I__3712\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18723\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__18728\,
            I => \N__18719\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__18723\,
            I => \N__18714\
        );

    \I__3709\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18711\
        );

    \I__3708\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18708\
        );

    \I__3707\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18703\
        );

    \I__3706\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18703\
        );

    \I__3705\ : Span4Mux_s3_v
    port map (
            O => \N__18714\,
            I => \N__18700\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__18711\,
            I => \sb_translator_1.num_ledsZ0Z_8\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__18708\,
            I => \sb_translator_1.num_ledsZ0Z_8\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__18703\,
            I => \sb_translator_1.num_ledsZ0Z_8\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__18700\,
            I => \sb_translator_1.num_ledsZ0Z_8\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__18691\,
            I => \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__18688\,
            I => \sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__18685\,
            I => \N__18677\
        );

    \I__3697\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18668\
        );

    \I__3696\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18668\
        );

    \I__3695\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18668\
        );

    \I__3694\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18668\
        );

    \I__3693\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18663\
        );

    \I__3692\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18663\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__18668\,
            I => \N__18660\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__18663\,
            I => \sb_translator_1.num_ledsZ0Z_3\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__18660\,
            I => \sb_translator_1.num_ledsZ0Z_3\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18652\
        );

    \I__3687\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18644\
        );

    \I__3686\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18644\
        );

    \I__3685\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18638\
        );

    \I__3684\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18638\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18635\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__18643\,
            I => \N__18631\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18626\
        );

    \I__3680\ : Span4Mux_s2_v
    port map (
            O => \N__18635\,
            I => \N__18626\
        );

    \I__3679\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18621\
        );

    \I__3678\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18621\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__18626\,
            I => \sb_translator_1.num_ledsZ0Z_4\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__18621\,
            I => \sb_translator_1.num_ledsZ0Z_4\
        );

    \I__3675\ : InMux
    port map (
            O => \N__18616\,
            I => \N__18613\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__18613\,
            I => \spi_slave_1.miso_data_outZ0Z_12\
        );

    \I__3673\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__18607\,
            I => \spi_slave_1.miso_data_outZ0Z_11\
        );

    \I__3671\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__18598\,
            I => \spi_slave_1.miso_RNOZ0Z_6\
        );

    \I__3668\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__18592\,
            I => \spi_slave_1.miso_data_outZ0Z_16\
        );

    \I__3666\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18586\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__18586\,
            I => \spi_slave_1.miso_data_outZ0Z_0\
        );

    \I__3664\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18575\
        );

    \I__3663\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18575\
        );

    \I__3662\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18572\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__18580\,
            I => \N__18568\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__18575\,
            I => \N__18565\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18560\
        );

    \I__3658\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18557\
        );

    \I__3657\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18554\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__18565\,
            I => \N__18551\
        );

    \I__3655\ : InMux
    port map (
            O => \N__18564\,
            I => \N__18546\
        );

    \I__3654\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18546\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__18560\,
            I => \N__18541\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18541\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__18554\,
            I => \spi_slave_1.bitcnt_txZ0Z_4\
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__18551\,
            I => \spi_slave_1.bitcnt_txZ0Z_4\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__18546\,
            I => \spi_slave_1.bitcnt_txZ0Z_4\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__18541\,
            I => \spi_slave_1.bitcnt_txZ0Z_4\
        );

    \I__3647\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18523\
        );

    \I__3646\ : InMux
    port map (
            O => \N__18531\,
            I => \N__18523\
        );

    \I__3645\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18523\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__18523\,
            I => \N__18518\
        );

    \I__3643\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18513\
        );

    \I__3642\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18513\
        );

    \I__3641\ : Span4Mux_h
    port map (
            O => \N__18518\,
            I => \N__18499\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18499\
        );

    \I__3639\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18496\
        );

    \I__3638\ : InMux
    port map (
            O => \N__18511\,
            I => \N__18493\
        );

    \I__3637\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18486\
        );

    \I__3636\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18486\
        );

    \I__3635\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18486\
        );

    \I__3634\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18477\
        );

    \I__3633\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18477\
        );

    \I__3632\ : InMux
    port map (
            O => \N__18505\,
            I => \N__18477\
        );

    \I__3631\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18477\
        );

    \I__3630\ : Span4Mux_h
    port map (
            O => \N__18499\,
            I => \N__18474\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__18496\,
            I => \spi_slave_1.bitcnt_txZ0Z_0\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__18493\,
            I => \spi_slave_1.bitcnt_txZ0Z_0\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__18486\,
            I => \spi_slave_1.bitcnt_txZ0Z_0\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__18477\,
            I => \spi_slave_1.bitcnt_txZ0Z_0\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__18474\,
            I => \spi_slave_1.bitcnt_txZ0Z_0\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__18463\,
            I => \spi_slave_1.N_58_0_cascade_\
        );

    \I__3623\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__18457\,
            I => \spi_slave_1.miso_data_outZ0Z_15\
        );

    \I__3621\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18451\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18448\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__18448\,
            I => \N__18445\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__18445\,
            I => \spi_slave_1.N_55_0\
        );

    \I__3617\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18439\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__18439\,
            I => \N__18435\
        );

    \I__3615\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18432\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__18435\,
            I => \spi_slave_1.mosi_data_inZ0Z_15\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__18432\,
            I => \spi_slave_1.mosi_data_inZ0Z_15\
        );

    \I__3612\ : CEMux
    port map (
            O => \N__18427\,
            I => \N__18415\
        );

    \I__3611\ : CEMux
    port map (
            O => \N__18426\,
            I => \N__18415\
        );

    \I__3610\ : CEMux
    port map (
            O => \N__18425\,
            I => \N__18415\
        );

    \I__3609\ : CEMux
    port map (
            O => \N__18424\,
            I => \N__18415\
        );

    \I__3608\ : GlobalMux
    port map (
            O => \N__18415\,
            I => \N__18412\
        );

    \I__3607\ : gio2CtrlBuf
    port map (
            O => \N__18412\,
            I => \spi_slave_1.un3_mosi_data_out_g\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_\
        );

    \I__3605\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18393\
        );

    \I__3604\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18393\
        );

    \I__3603\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18393\
        );

    \I__3602\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18393\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__18402\,
            I => \N__18389\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__18393\,
            I => \N__18386\
        );

    \I__3599\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18381\
        );

    \I__3598\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18381\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__18386\,
            I => \sb_translator_1.num_ledsZ0Z_5\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__18381\,
            I => \sb_translator_1.num_ledsZ0Z_5\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_\
        );

    \I__3594\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18368\
        );

    \I__3593\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18363\
        );

    \I__3592\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18363\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__18368\,
            I => \demux.N_239\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__18363\,
            I => \demux.N_239\
        );

    \I__3589\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18353\
        );

    \I__3588\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18348\
        );

    \I__3587\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18348\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__18353\,
            I => \demux.N_241\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__18348\,
            I => \demux.N_241\
        );

    \I__3584\ : InMux
    port map (
            O => \N__18343\,
            I => \N__18336\
        );

    \I__3583\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18336\
        );

    \I__3582\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18333\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__18336\,
            I => \demux.N_915\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__18333\,
            I => \demux.N_915\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__3578\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18317\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18317\
        );

    \I__3576\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18312\
        );

    \I__3575\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18312\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__18317\,
            I => ram_sel_12
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__18312\,
            I => ram_sel_12
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__18307\,
            I => \demux.N_915_cascade_\
        );

    \I__3571\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18296\
        );

    \I__3570\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18296\
        );

    \I__3569\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18291\
        );

    \I__3568\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18291\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__18296\,
            I => ram_sel_2
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__18291\,
            I => ram_sel_2
        );

    \I__3565\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18281\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__18285\,
            I => \N__18278\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__18284\,
            I => \N__18275\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__18281\,
            I => \N__18270\
        );

    \I__3561\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18263\
        );

    \I__3560\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18263\
        );

    \I__3559\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18263\
        );

    \I__3558\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18260\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__18270\,
            I => ram_sel_3
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__18263\,
            I => ram_sel_3
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__18260\,
            I => ram_sel_3
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__18253\,
            I => \N__18247\
        );

    \I__3553\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18239\
        );

    \I__3552\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18239\
        );

    \I__3551\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18239\
        );

    \I__3550\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18234\
        );

    \I__3549\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18234\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__18239\,
            I => ram_sel_8
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__18234\,
            I => ram_sel_8
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__18228\,
            I => \N__18220\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__18227\,
            I => \N__18217\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__18226\,
            I => \N__18214\
        );

    \I__3542\ : CascadeBuf
    port map (
            O => \N__18223\,
            I => \N__18211\
        );

    \I__3541\ : CascadeBuf
    port map (
            O => \N__18220\,
            I => \N__18208\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__18217\,
            I => \N__18205\
        );

    \I__3539\ : CascadeBuf
    port map (
            O => \N__18214\,
            I => \N__18202\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__18211\,
            I => \N__18199\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__18208\,
            I => \N__18196\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__18205\,
            I => \N__18193\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__18202\,
            I => \N__18190\
        );

    \I__3534\ : CascadeBuf
    port map (
            O => \N__18199\,
            I => \N__18187\
        );

    \I__3533\ : CascadeBuf
    port map (
            O => \N__18196\,
            I => \N__18184\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__18193\,
            I => \N__18181\
        );

    \I__3531\ : CascadeBuf
    port map (
            O => \N__18190\,
            I => \N__18178\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__18187\,
            I => \N__18175\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__18184\,
            I => \N__18172\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__18181\,
            I => \N__18169\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__18178\,
            I => \N__18166\
        );

    \I__3526\ : CascadeBuf
    port map (
            O => \N__18175\,
            I => \N__18163\
        );

    \I__3525\ : CascadeBuf
    port map (
            O => \N__18172\,
            I => \N__18160\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__18169\,
            I => \N__18157\
        );

    \I__3523\ : CascadeBuf
    port map (
            O => \N__18166\,
            I => \N__18154\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__18163\,
            I => \N__18151\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__18160\,
            I => \N__18148\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__18157\,
            I => \N__18145\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__18154\,
            I => \N__18142\
        );

    \I__3518\ : CascadeBuf
    port map (
            O => \N__18151\,
            I => \N__18139\
        );

    \I__3517\ : CascadeBuf
    port map (
            O => \N__18148\,
            I => \N__18136\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__18145\,
            I => \N__18133\
        );

    \I__3515\ : CascadeBuf
    port map (
            O => \N__18142\,
            I => \N__18130\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__18139\,
            I => \N__18127\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__18136\,
            I => \N__18124\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__18133\,
            I => \N__18121\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__18130\,
            I => \N__18118\
        );

    \I__3510\ : CascadeBuf
    port map (
            O => \N__18127\,
            I => \N__18115\
        );

    \I__3509\ : CascadeBuf
    port map (
            O => \N__18124\,
            I => \N__18112\
        );

    \I__3508\ : CascadeBuf
    port map (
            O => \N__18121\,
            I => \N__18109\
        );

    \I__3507\ : CascadeBuf
    port map (
            O => \N__18118\,
            I => \N__18106\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18103\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \N__18100\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__18109\,
            I => \N__18097\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18094\
        );

    \I__3502\ : CascadeBuf
    port map (
            O => \N__18103\,
            I => \N__18091\
        );

    \I__3501\ : CascadeBuf
    port map (
            O => \N__18100\,
            I => \N__18088\
        );

    \I__3500\ : CascadeBuf
    port map (
            O => \N__18097\,
            I => \N__18085\
        );

    \I__3499\ : CascadeBuf
    port map (
            O => \N__18094\,
            I => \N__18082\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__18091\,
            I => \N__18079\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__18088\,
            I => \N__18076\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__18085\,
            I => \N__18073\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__18082\,
            I => \N__18070\
        );

    \I__3494\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18067\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18064\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18061\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18058\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18067\,
            I => \N__18052\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__18064\,
            I => \N__18052\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__18061\,
            I => \N__18047\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__18058\,
            I => \N__18047\
        );

    \I__3486\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18044\
        );

    \I__3485\ : Span4Mux_s2_v
    port map (
            O => \N__18052\,
            I => \N__18041\
        );

    \I__3484\ : Span4Mux_s2_v
    port map (
            O => \N__18047\,
            I => \N__18038\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__18044\,
            I => addr_out_8
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__18041\,
            I => addr_out_8
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__18038\,
            I => addr_out_8
        );

    \I__3480\ : CEMux
    port map (
            O => \N__18031\,
            I => \N__18028\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__18028\,
            I => \N__18024\
        );

    \I__3478\ : CEMux
    port map (
            O => \N__18027\,
            I => \N__18021\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__18024\,
            I => \N__18018\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__18021\,
            I => \N__18015\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__18018\,
            I => \sb_translator_1.state_RNI88IGAZ0Z_0\
        );

    \I__3474\ : Odrv12
    port map (
            O => \N__18015\,
            I => \sb_translator_1.state_RNI88IGAZ0Z_0\
        );

    \I__3473\ : IoInMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__18004\
        );

    \I__3471\ : Span4Mux_s0_v
    port map (
            O => \N__18004\,
            I => \N__18001\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__18001\,
            I => \sb_translator_1.state_leds_2_sqmuxa\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__17998\,
            I => \N__17994\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__17997\,
            I => \N__17990\
        );

    \I__3467\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17985\
        );

    \I__3466\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17985\
        );

    \I__3465\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17982\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__17985\,
            I => \N__17979\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__17982\,
            I => \sb_translator_1.state_ledsZ0\
        );

    \I__3462\ : Odrv12
    port map (
            O => \N__17979\,
            I => \sb_translator_1.state_ledsZ0\
        );

    \I__3461\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17971\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__17971\,
            I => \spi_slave_1.miso_data_outZ0Z_9\
        );

    \I__3459\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__17965\,
            I => \spi_slave_1.miso_data_outZ0Z_10\
        );

    \I__3457\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17959\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__17959\,
            I => \N__17956\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__17956\,
            I => \spi_slave_1.miso_RNOZ0Z_13\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__17953\,
            I => \demux.N_242_cascade_\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__17950\,
            I => \demux.N_424_i_0_a2Z0Z_34_cascade_\
        );

    \I__3452\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17938\
        );

    \I__3451\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17938\
        );

    \I__3450\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17928\
        );

    \I__3449\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17928\
        );

    \I__3448\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17928\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17925\
        );

    \I__3446\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17918\
        );

    \I__3445\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17918\
        );

    \I__3444\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17918\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__17928\,
            I => \N__17915\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__17925\,
            I => \N__17912\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__17918\,
            I => \demux.N_424_i_0_aZ0Z2\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__17915\,
            I => \demux.N_424_i_0_aZ0Z2\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__17912\,
            I => \demux.N_424_i_0_aZ0Z2\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17901\
        );

    \I__3437\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17898\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__17901\,
            I => \demux.N_242\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__17898\,
            I => \demux.N_242\
        );

    \I__3434\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17884\
        );

    \I__3433\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17884\
        );

    \I__3432\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17884\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__17884\,
            I => \demux.N_916\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__17881\,
            I => \N__17876\
        );

    \I__3429\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17872\
        );

    \I__3428\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17865\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17865\
        );

    \I__3426\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17865\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__17872\,
            I => ram_sel_5
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__17865\,
            I => ram_sel_5
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__17860\,
            I => \demux.N_916_cascade_\
        );

    \I__3422\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17851\
        );

    \I__3421\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17848\
        );

    \I__3420\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17843\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17843\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__17851\,
            I => ram_sel_1
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__17848\,
            I => ram_sel_1
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__17843\,
            I => ram_sel_1
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__17836\,
            I => \sb_translator_1.num_leds_1_sqmuxa_cascade_\
        );

    \I__3414\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17826\
        );

    \I__3413\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17826\
        );

    \I__3412\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17823\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__17826\,
            I => \N__17818\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__17823\,
            I => \N__17818\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__17818\,
            I => \N__17815\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__17815\,
            I => \sb_translator_1.send_leds_n_1_sqmuxa\
        );

    \I__3407\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17809\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__17809\,
            I => \sb_translator_1.N_59\
        );

    \I__3405\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17803\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17800\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__17800\,
            I => \N__17797\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__17797\,
            I => miso_data_in_0
        );

    \I__3401\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17789\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \N__17785\
        );

    \I__3399\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17782\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17779\
        );

    \I__3397\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17774\
        );

    \I__3396\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17774\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__17782\,
            I => \N__17771\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__17779\,
            I => \N__17768\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__17774\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5\
        );

    \I__3392\ : Odrv4
    port map (
            O => \N__17771\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__17768\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5\
        );

    \I__3390\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17758\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17754\
        );

    \I__3388\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17751\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__17754\,
            I => \N__17746\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__17751\,
            I => \N__17743\
        );

    \I__3385\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17740\
        );

    \I__3384\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17737\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__17746\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__17743\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__17740\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__17737\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__17728\,
            I => \N__17724\
        );

    \I__3378\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17721\
        );

    \I__3377\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17716\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__17721\,
            I => \N__17713\
        );

    \I__3375\ : InMux
    port map (
            O => \N__17720\,
            I => \N__17708\
        );

    \I__3374\ : InMux
    port map (
            O => \N__17719\,
            I => \N__17708\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__17716\,
            I => \N__17705\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__17713\,
            I => \N__17702\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__17708\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__17705\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__17702\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0\
        );

    \I__3368\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17683\
        );

    \I__3367\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17683\
        );

    \I__3366\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17683\
        );

    \I__3365\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17683\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__17683\,
            I => \N__17676\
        );

    \I__3363\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17671\
        );

    \I__3362\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17671\
        );

    \I__3361\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17668\
        );

    \I__3360\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17665\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__17676\,
            I => \N__17660\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17660\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17655\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17655\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__17660\,
            I => \N__17652\
        );

    \I__3354\ : Span4Mux_v
    port map (
            O => \N__17655\,
            I => \N__17649\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__17652\,
            I => mosi_data_out_18
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__17649\,
            I => mosi_data_out_18
        );

    \I__3351\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17636\
        );

    \I__3350\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17636\
        );

    \I__3349\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17631\
        );

    \I__3348\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17631\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17624\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__17631\,
            I => \N__17624\
        );

    \I__3345\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17617\
        );

    \I__3344\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17617\
        );

    \I__3343\ : Span4Mux_v
    port map (
            O => \N__17624\,
            I => \N__17614\
        );

    \I__3342\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17609\
        );

    \I__3341\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17609\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17606\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__17614\,
            I => \N__17601\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__17609\,
            I => \N__17601\
        );

    \I__3337\ : Span12Mux_s11_h
    port map (
            O => \N__17606\,
            I => \N__17598\
        );

    \I__3336\ : Span4Mux_v
    port map (
            O => \N__17601\,
            I => \N__17595\
        );

    \I__3335\ : Odrv12
    port map (
            O => \N__17598\,
            I => mosi_data_out_19
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__17595\,
            I => mosi_data_out_19
        );

    \I__3333\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17578\
        );

    \I__3332\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17578\
        );

    \I__3331\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17578\
        );

    \I__3330\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17578\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17573\
        );

    \I__3328\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17568\
        );

    \I__3327\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17565\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__17573\,
            I => \N__17562\
        );

    \I__3325\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17557\
        );

    \I__3324\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17557\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__17568\,
            I => \N__17552\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__17565\,
            I => \N__17552\
        );

    \I__3321\ : Span4Mux_h
    port map (
            O => \N__17562\,
            I => \N__17547\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__17557\,
            I => \N__17547\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__17552\,
            I => \N__17544\
        );

    \I__3318\ : Span4Mux_v
    port map (
            O => \N__17547\,
            I => \N__17541\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__17544\,
            I => mosi_data_out_20
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__17541\,
            I => mosi_data_out_20
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__17536\,
            I => \N__17533\
        );

    \I__3314\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17530\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__17530\,
            I => \N__17524\
        );

    \I__3312\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17521\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__17528\,
            I => \N__17518\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__17527\,
            I => \N__17515\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__17524\,
            I => \N__17512\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__17521\,
            I => \N__17509\
        );

    \I__3307\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17504\
        );

    \I__3306\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17504\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__17512\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__17509\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__17504\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \demux.N_238_cascade_\
        );

    \I__3301\ : CEMux
    port map (
            O => \N__17494\,
            I => \N__17490\
        );

    \I__3300\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17487\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17484\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__17487\,
            I => \N__17479\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__17484\,
            I => \N__17476\
        );

    \I__3296\ : CEMux
    port map (
            O => \N__17483\,
            I => \N__17473\
        );

    \I__3295\ : CEMux
    port map (
            O => \N__17482\,
            I => \N__17470\
        );

    \I__3294\ : Span12Mux_s9_h
    port map (
            O => \N__17479\,
            I => \N__17467\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__17476\,
            I => \sb_translator_1.N_58\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__17473\,
            I => \sb_translator_1.N_58\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__17470\,
            I => \sb_translator_1.N_58\
        );

    \I__3290\ : Odrv12
    port map (
            O => \N__17467\,
            I => \sb_translator_1.N_58\
        );

    \I__3289\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17455\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__17455\,
            I => \sb_translator_1.state_RNIEL0N9_0Z0Z_6\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__17452\,
            I => \N__17444\
        );

    \I__3286\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17432\
        );

    \I__3285\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17432\
        );

    \I__3284\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17432\
        );

    \I__3283\ : InMux
    port map (
            O => \N__17448\,
            I => \N__17432\
        );

    \I__3282\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17432\
        );

    \I__3281\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17427\
        );

    \I__3280\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17427\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17424\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__17427\,
            I => \sb_translator_1.cnt_ram_readZ0Z_0\
        );

    \I__3277\ : Odrv12
    port map (
            O => \N__17424\,
            I => \sb_translator_1.cnt_ram_readZ0Z_0\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__17418\,
            I => \N__17410\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \N__17407\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__17416\,
            I => \N__17403\
        );

    \I__3272\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17399\
        );

    \I__3271\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17388\
        );

    \I__3270\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17388\
        );

    \I__3269\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17388\
        );

    \I__3268\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17388\
        );

    \I__3267\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17388\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17383\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__17388\,
            I => \N__17383\
        );

    \I__3264\ : Odrv12
    port map (
            O => \N__17383\,
            I => \sb_translator_1.cnt_ram_readZ0Z_1\
        );

    \I__3263\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__17377\,
            I => \N__17374\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__17371\,
            I => demux_data_in_42
        );

    \I__3259\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17364\
        );

    \I__3258\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17361\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__17364\,
            I => \N__17355\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__17361\,
            I => \N__17352\
        );

    \I__3255\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17347\
        );

    \I__3254\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17347\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17343\
        );

    \I__3252\ : Span4Mux_v
    port map (
            O => \N__17355\,
            I => \N__17338\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__17352\,
            I => \N__17338\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__17347\,
            I => \N__17335\
        );

    \I__3249\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17332\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17329\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__17338\,
            I => \sb_translator_1.cntZ0Z_11\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__17335\,
            I => \sb_translator_1.cntZ0Z_11\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__17332\,
            I => \sb_translator_1.cntZ0Z_11\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__17329\,
            I => \sb_translator_1.cntZ0Z_11\
        );

    \I__3243\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17316\
        );

    \I__3242\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17313\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17308\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__17313\,
            I => \N__17305\
        );

    \I__3239\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17300\
        );

    \I__3238\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17300\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__17308\,
            I => \N__17293\
        );

    \I__3236\ : Span4Mux_v
    port map (
            O => \N__17305\,
            I => \N__17293\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__17300\,
            I => \N__17293\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__17293\,
            I => \N__17288\
        );

    \I__3233\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17285\
        );

    \I__3232\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17282\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__17288\,
            I => \sb_translator_1.cntZ0Z_10\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__17285\,
            I => \sb_translator_1.cntZ0Z_10\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__17282\,
            I => \sb_translator_1.cntZ0Z_10\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__17275\,
            I => \N__17272\
        );

    \I__3227\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17269\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17266\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__17266\,
            I => \N__17262\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__17265\,
            I => \N__17259\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__17262\,
            I => \N__17256\
        );

    \I__3222\ : InMux
    port map (
            O => \N__17259\,
            I => \N__17253\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__17256\,
            I => \sb_translator_1.ram_we_6_0_0_a2_0_6\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__17253\,
            I => \sb_translator_1.ram_we_6_0_0_a2_0_6\
        );

    \I__3219\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17245\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17242\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__17242\,
            I => \N__17239\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__17239\,
            I => miso_data_in_2
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__17236\,
            I => \N__17229\
        );

    \I__3214\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17224\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__17234\,
            I => \N__17217\
        );

    \I__3212\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17210\
        );

    \I__3211\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17210\
        );

    \I__3210\ : InMux
    port map (
            O => \N__17229\,
            I => \N__17210\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \N__17207\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__17227\,
            I => \N__17204\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__17224\,
            I => \N__17193\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__17223\,
            I => \N__17190\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__17222\,
            I => \N__17187\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__17221\,
            I => \N__17184\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__17220\,
            I => \N__17181\
        );

    \I__3202\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17174\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__17210\,
            I => \N__17171\
        );

    \I__3200\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17164\
        );

    \I__3199\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17164\
        );

    \I__3198\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17164\
        );

    \I__3197\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17149\
        );

    \I__3196\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17149\
        );

    \I__3195\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17149\
        );

    \I__3194\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17149\
        );

    \I__3193\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17149\
        );

    \I__3192\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17149\
        );

    \I__3191\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17149\
        );

    \I__3190\ : Span4Mux_v
    port map (
            O => \N__17193\,
            I => \N__17146\
        );

    \I__3189\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17129\
        );

    \I__3188\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17129\
        );

    \I__3187\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17129\
        );

    \I__3186\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17129\
        );

    \I__3185\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17129\
        );

    \I__3184\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17129\
        );

    \I__3183\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17129\
        );

    \I__3182\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17129\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__17174\,
            I => \N__17126\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__17171\,
            I => \N__17123\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__17164\,
            I => \N__17116\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__17149\,
            I => \N__17116\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__17146\,
            I => \N__17116\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__17129\,
            I => mosi_data_out_22
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__17126\,
            I => mosi_data_out_22
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__17123\,
            I => mosi_data_out_22
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__17116\,
            I => mosi_data_out_22
        );

    \I__3172\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17083\
        );

    \I__3171\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17083\
        );

    \I__3170\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17083\
        );

    \I__3169\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17068\
        );

    \I__3168\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17068\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17068\
        );

    \I__3166\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17068\
        );

    \I__3165\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17068\
        );

    \I__3164\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17068\
        );

    \I__3163\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17068\
        );

    \I__3162\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17051\
        );

    \I__3161\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17051\
        );

    \I__3160\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17051\
        );

    \I__3159\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17051\
        );

    \I__3158\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17051\
        );

    \I__3157\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17051\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17051\
        );

    \I__3155\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17051\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__17083\,
            I => \N__17043\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17043\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__17051\,
            I => \N__17043\
        );

    \I__3151\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17040\
        );

    \I__3150\ : Span4Mux_v
    port map (
            O => \N__17043\,
            I => \N__17037\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17034\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__17037\,
            I => \sb_translator_1.N_1087\
        );

    \I__3147\ : Odrv12
    port map (
            O => \N__17034\,
            I => \sb_translator_1.N_1087\
        );

    \I__3146\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17026\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__17026\,
            I => \N__17021\
        );

    \I__3144\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17018\
        );

    \I__3143\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17015\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__17021\,
            I => mosi_data_out_3
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__17018\,
            I => mosi_data_out_3
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__17015\,
            I => mosi_data_out_3
        );

    \I__3139\ : InMux
    port map (
            O => \N__17008\,
            I => \N__17005\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__17005\,
            I => \sb_translator_1.instr_tmpZ1Z_3\
        );

    \I__3137\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16997\
        );

    \I__3136\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16994\
        );

    \I__3135\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16991\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16988\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__16994\,
            I => mosi_data_out_4
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__16991\,
            I => mosi_data_out_4
        );

    \I__3131\ : Odrv12
    port map (
            O => \N__16988\,
            I => mosi_data_out_4
        );

    \I__3130\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16978\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__16978\,
            I => \sb_translator_1.instr_tmpZ1Z_4\
        );

    \I__3128\ : CEMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__16972\,
            I => \N__16968\
        );

    \I__3126\ : CEMux
    port map (
            O => \N__16971\,
            I => \N__16965\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__16968\,
            I => \N__16960\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__16965\,
            I => \N__16960\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__16960\,
            I => \N__16957\
        );

    \I__3122\ : Span4Mux_s1_h
    port map (
            O => \N__16957\,
            I => \N__16954\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__16954\,
            I => \sb_translator_1.state_RNIKJOCZ0Z_5\
        );

    \I__3120\ : InMux
    port map (
            O => \N__16951\,
            I => \N__16947\
        );

    \I__3119\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16942\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__16947\,
            I => \N__16939\
        );

    \I__3117\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16936\
        );

    \I__3116\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16933\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__16942\,
            I => \N__16930\
        );

    \I__3114\ : Span4Mux_h
    port map (
            O => \N__16939\,
            I => \N__16927\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__16936\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__16933\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\
        );

    \I__3111\ : Odrv12
    port map (
            O => \N__16930\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__16927\,
            I => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__16918\,
            I => \N__16912\
        );

    \I__3108\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16907\
        );

    \I__3107\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16907\
        );

    \I__3106\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16904\
        );

    \I__3105\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16901\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16898\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16895\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__16901\,
            I => \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11\
        );

    \I__3101\ : Odrv4
    port map (
            O => \N__16898\,
            I => \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__16895\,
            I => \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11\
        );

    \I__3099\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__16885\,
            I => \N__16882\
        );

    \I__3097\ : Span4Mux_v
    port map (
            O => \N__16882\,
            I => \N__16878\
        );

    \I__3096\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16875\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__16875\,
            I => \sb_translator_1.cnt19_cry_18_THRU_CO\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__16872\,
            I => \sb_translator_1.cnt19_cry_18_THRU_CO\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__16867\,
            I => \sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_\
        );

    \I__3091\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16857\
        );

    \I__3090\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16854\
        );

    \I__3089\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16845\
        );

    \I__3088\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16845\
        );

    \I__3087\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16845\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__16857\,
            I => \N__16837\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__16854\,
            I => \N__16837\
        );

    \I__3084\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16834\
        );

    \I__3083\ : InMux
    port map (
            O => \N__16852\,
            I => \N__16831\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__16845\,
            I => \N__16828\
        );

    \I__3081\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16818\
        );

    \I__3080\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16818\
        );

    \I__3079\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16818\
        );

    \I__3078\ : Span12Mux_h
    port map (
            O => \N__16837\,
            I => \N__16815\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__16834\,
            I => \N__16812\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__16831\,
            I => \N__16807\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__16828\,
            I => \N__16807\
        );

    \I__3074\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16800\
        );

    \I__3073\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16800\
        );

    \I__3072\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16800\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__16818\,
            I => mosi_rx
        );

    \I__3070\ : Odrv12
    port map (
            O => \N__16815\,
            I => mosi_rx
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__16812\,
            I => mosi_rx
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__16807\,
            I => mosi_rx
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__16800\,
            I => mosi_rx
        );

    \I__3066\ : CEMux
    port map (
            O => \N__16789\,
            I => \N__16786\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16781\
        );

    \I__3064\ : CEMux
    port map (
            O => \N__16785\,
            I => \N__16778\
        );

    \I__3063\ : CEMux
    port map (
            O => \N__16784\,
            I => \N__16775\
        );

    \I__3062\ : Span4Mux_h
    port map (
            O => \N__16781\,
            I => \N__16772\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__16778\,
            I => \N__16769\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16766\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__16772\,
            I => \sb_translator_1.state_RNIOH7V9Z0Z_0\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__16769\,
            I => \sb_translator_1.state_RNIOH7V9Z0Z_0\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__16766\,
            I => \sb_translator_1.state_RNIOH7V9Z0Z_0\
        );

    \I__3056\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16756\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__16756\,
            I => \N__16753\
        );

    \I__3054\ : Odrv12
    port map (
            O => \N__16753\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_5\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__16750\,
            I => \N__16747\
        );

    \I__3052\ : CascadeBuf
    port map (
            O => \N__16747\,
            I => \N__16744\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__16744\,
            I => \N__16739\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__16743\,
            I => \N__16736\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__16742\,
            I => \N__16733\
        );

    \I__3048\ : CascadeBuf
    port map (
            O => \N__16739\,
            I => \N__16730\
        );

    \I__3047\ : CascadeBuf
    port map (
            O => \N__16736\,
            I => \N__16727\
        );

    \I__3046\ : CascadeBuf
    port map (
            O => \N__16733\,
            I => \N__16723\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__16730\,
            I => \N__16720\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \N__16717\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__16726\,
            I => \N__16714\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__16723\,
            I => \N__16711\
        );

    \I__3041\ : CascadeBuf
    port map (
            O => \N__16720\,
            I => \N__16708\
        );

    \I__3040\ : CascadeBuf
    port map (
            O => \N__16717\,
            I => \N__16705\
        );

    \I__3039\ : CascadeBuf
    port map (
            O => \N__16714\,
            I => \N__16702\
        );

    \I__3038\ : CascadeBuf
    port map (
            O => \N__16711\,
            I => \N__16699\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__16708\,
            I => \N__16696\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__16705\,
            I => \N__16693\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__16702\,
            I => \N__16690\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__16699\,
            I => \N__16687\
        );

    \I__3033\ : CascadeBuf
    port map (
            O => \N__16696\,
            I => \N__16684\
        );

    \I__3032\ : CascadeBuf
    port map (
            O => \N__16693\,
            I => \N__16681\
        );

    \I__3031\ : CascadeBuf
    port map (
            O => \N__16690\,
            I => \N__16678\
        );

    \I__3030\ : CascadeBuf
    port map (
            O => \N__16687\,
            I => \N__16675\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__16684\,
            I => \N__16672\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__16681\,
            I => \N__16669\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \N__16666\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__16675\,
            I => \N__16663\
        );

    \I__3025\ : CascadeBuf
    port map (
            O => \N__16672\,
            I => \N__16660\
        );

    \I__3024\ : CascadeBuf
    port map (
            O => \N__16669\,
            I => \N__16657\
        );

    \I__3023\ : CascadeBuf
    port map (
            O => \N__16666\,
            I => \N__16654\
        );

    \I__3022\ : CascadeBuf
    port map (
            O => \N__16663\,
            I => \N__16651\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__16660\,
            I => \N__16648\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__16657\,
            I => \N__16645\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__16654\,
            I => \N__16642\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__16651\,
            I => \N__16639\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__16648\,
            I => \N__16636\
        );

    \I__3016\ : CascadeBuf
    port map (
            O => \N__16645\,
            I => \N__16633\
        );

    \I__3015\ : CascadeBuf
    port map (
            O => \N__16642\,
            I => \N__16630\
        );

    \I__3014\ : CascadeBuf
    port map (
            O => \N__16639\,
            I => \N__16627\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__16636\,
            I => \N__16624\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__16633\,
            I => \N__16621\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__16630\,
            I => \N__16618\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__16627\,
            I => \N__16615\
        );

    \I__3009\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16612\
        );

    \I__3008\ : CascadeBuf
    port map (
            O => \N__16621\,
            I => \N__16609\
        );

    \I__3007\ : CascadeBuf
    port map (
            O => \N__16618\,
            I => \N__16606\
        );

    \I__3006\ : CascadeBuf
    port map (
            O => \N__16615\,
            I => \N__16603\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16600\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__16609\,
            I => \N__16597\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__16606\,
            I => \N__16594\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__16603\,
            I => \N__16591\
        );

    \I__3001\ : Span4Mux_s1_v
    port map (
            O => \N__16600\,
            I => \N__16587\
        );

    \I__3000\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16584\
        );

    \I__2999\ : CascadeBuf
    port map (
            O => \N__16594\,
            I => \N__16581\
        );

    \I__2998\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16578\
        );

    \I__2997\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16575\
        );

    \I__2996\ : Span4Mux_s2_h
    port map (
            O => \N__16587\,
            I => \N__16570\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__16584\,
            I => \N__16570\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__16581\,
            I => \N__16567\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16564\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16559\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__16570\,
            I => \N__16559\
        );

    \I__2990\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16556\
        );

    \I__2989\ : Span4Mux_s1_v
    port map (
            O => \N__16564\,
            I => \N__16549\
        );

    \I__2988\ : Span4Mux_h
    port map (
            O => \N__16559\,
            I => \N__16549\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__16556\,
            I => \N__16549\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__16549\,
            I => \N__16546\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__16546\,
            I => \N__16543\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__16543\,
            I => addr_out_5
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__16540\,
            I => \N__16535\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__16539\,
            I => \N__16532\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__16538\,
            I => \N__16529\
        );

    \I__2980\ : CascadeBuf
    port map (
            O => \N__16535\,
            I => \N__16526\
        );

    \I__2979\ : CascadeBuf
    port map (
            O => \N__16532\,
            I => \N__16522\
        );

    \I__2978\ : CascadeBuf
    port map (
            O => \N__16529\,
            I => \N__16519\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__16526\,
            I => \N__16516\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__16525\,
            I => \N__16513\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__16522\,
            I => \N__16510\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__16519\,
            I => \N__16507\
        );

    \I__2973\ : CascadeBuf
    port map (
            O => \N__16516\,
            I => \N__16504\
        );

    \I__2972\ : CascadeBuf
    port map (
            O => \N__16513\,
            I => \N__16501\
        );

    \I__2971\ : CascadeBuf
    port map (
            O => \N__16510\,
            I => \N__16498\
        );

    \I__2970\ : CascadeBuf
    port map (
            O => \N__16507\,
            I => \N__16495\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__16504\,
            I => \N__16492\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__16501\,
            I => \N__16489\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__16498\,
            I => \N__16486\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__16495\,
            I => \N__16483\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__16492\,
            I => \N__16480\
        );

    \I__2964\ : CascadeBuf
    port map (
            O => \N__16489\,
            I => \N__16477\
        );

    \I__2963\ : CascadeBuf
    port map (
            O => \N__16486\,
            I => \N__16474\
        );

    \I__2962\ : CascadeBuf
    port map (
            O => \N__16483\,
            I => \N__16471\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16468\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__16477\,
            I => \N__16465\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__16474\,
            I => \N__16462\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__16471\,
            I => \N__16459\
        );

    \I__2957\ : CascadeBuf
    port map (
            O => \N__16468\,
            I => \N__16456\
        );

    \I__2956\ : CascadeBuf
    port map (
            O => \N__16465\,
            I => \N__16453\
        );

    \I__2955\ : CascadeBuf
    port map (
            O => \N__16462\,
            I => \N__16450\
        );

    \I__2954\ : CascadeBuf
    port map (
            O => \N__16459\,
            I => \N__16447\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__16456\,
            I => \N__16444\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__16453\,
            I => \N__16441\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \N__16438\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__16447\,
            I => \N__16435\
        );

    \I__2949\ : CascadeBuf
    port map (
            O => \N__16444\,
            I => \N__16432\
        );

    \I__2948\ : CascadeBuf
    port map (
            O => \N__16441\,
            I => \N__16429\
        );

    \I__2947\ : CascadeBuf
    port map (
            O => \N__16438\,
            I => \N__16426\
        );

    \I__2946\ : CascadeBuf
    port map (
            O => \N__16435\,
            I => \N__16423\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__16432\,
            I => \N__16420\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__16429\,
            I => \N__16417\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__16426\,
            I => \N__16414\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__16423\,
            I => \N__16411\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__16420\,
            I => \N__16408\
        );

    \I__2940\ : CascadeBuf
    port map (
            O => \N__16417\,
            I => \N__16405\
        );

    \I__2939\ : CascadeBuf
    port map (
            O => \N__16414\,
            I => \N__16402\
        );

    \I__2938\ : CascadeBuf
    port map (
            O => \N__16411\,
            I => \N__16399\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__16408\,
            I => \N__16396\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \N__16393\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16390\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__16399\,
            I => \N__16387\
        );

    \I__2933\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16383\
        );

    \I__2932\ : CascadeBuf
    port map (
            O => \N__16393\,
            I => \N__16380\
        );

    \I__2931\ : InMux
    port map (
            O => \N__16390\,
            I => \N__16377\
        );

    \I__2930\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16374\
        );

    \I__2929\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16371\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__16383\,
            I => \N__16368\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__16380\,
            I => \N__16365\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__16377\,
            I => \N__16362\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__16374\,
            I => \N__16359\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__16371\,
            I => \N__16354\
        );

    \I__2923\ : Span4Mux_h
    port map (
            O => \N__16368\,
            I => \N__16354\
        );

    \I__2922\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16351\
        );

    \I__2921\ : Span4Mux_s3_v
    port map (
            O => \N__16362\,
            I => \N__16348\
        );

    \I__2920\ : Span4Mux_s1_v
    port map (
            O => \N__16359\,
            I => \N__16341\
        );

    \I__2919\ : Span4Mux_h
    port map (
            O => \N__16354\,
            I => \N__16341\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__16351\,
            I => \N__16341\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__16348\,
            I => \N__16338\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__16341\,
            I => \N__16335\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__16338\,
            I => \N__16332\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__16335\,
            I => \N__16329\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__16332\,
            I => addr_out_6
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__16329\,
            I => addr_out_6
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__16324\,
            I => \N__16319\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__16323\,
            I => \N__16316\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__16322\,
            I => \N__16313\
        );

    \I__2908\ : CascadeBuf
    port map (
            O => \N__16319\,
            I => \N__16310\
        );

    \I__2907\ : CascadeBuf
    port map (
            O => \N__16316\,
            I => \N__16306\
        );

    \I__2906\ : CascadeBuf
    port map (
            O => \N__16313\,
            I => \N__16303\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N__16300\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16297\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__16306\,
            I => \N__16294\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__16303\,
            I => \N__16291\
        );

    \I__2901\ : CascadeBuf
    port map (
            O => \N__16300\,
            I => \N__16288\
        );

    \I__2900\ : CascadeBuf
    port map (
            O => \N__16297\,
            I => \N__16285\
        );

    \I__2899\ : CascadeBuf
    port map (
            O => \N__16294\,
            I => \N__16282\
        );

    \I__2898\ : CascadeBuf
    port map (
            O => \N__16291\,
            I => \N__16279\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__16288\,
            I => \N__16276\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__16285\,
            I => \N__16273\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__16282\,
            I => \N__16270\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__16279\,
            I => \N__16267\
        );

    \I__2893\ : CascadeBuf
    port map (
            O => \N__16276\,
            I => \N__16264\
        );

    \I__2892\ : CascadeBuf
    port map (
            O => \N__16273\,
            I => \N__16261\
        );

    \I__2891\ : CascadeBuf
    port map (
            O => \N__16270\,
            I => \N__16258\
        );

    \I__2890\ : CascadeBuf
    port map (
            O => \N__16267\,
            I => \N__16255\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__16264\,
            I => \N__16252\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__16261\,
            I => \N__16249\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__16258\,
            I => \N__16246\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__16255\,
            I => \N__16243\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__16252\,
            I => \N__16240\
        );

    \I__2884\ : CascadeBuf
    port map (
            O => \N__16249\,
            I => \N__16237\
        );

    \I__2883\ : CascadeBuf
    port map (
            O => \N__16246\,
            I => \N__16234\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__16243\,
            I => \N__16231\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__16240\,
            I => \N__16228\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16225\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__16234\,
            I => \N__16222\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__16231\,
            I => \N__16219\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__16228\,
            I => \N__16216\
        );

    \I__2876\ : CascadeBuf
    port map (
            O => \N__16225\,
            I => \N__16213\
        );

    \I__2875\ : CascadeBuf
    port map (
            O => \N__16222\,
            I => \N__16210\
        );

    \I__2874\ : CascadeBuf
    port map (
            O => \N__16219\,
            I => \N__16207\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__16216\,
            I => \N__16204\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16201\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__16210\,
            I => \N__16198\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__16207\,
            I => \N__16195\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__16204\,
            I => \N__16192\
        );

    \I__2868\ : CascadeBuf
    port map (
            O => \N__16201\,
            I => \N__16189\
        );

    \I__2867\ : CascadeBuf
    port map (
            O => \N__16198\,
            I => \N__16186\
        );

    \I__2866\ : CascadeBuf
    port map (
            O => \N__16195\,
            I => \N__16183\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__16192\,
            I => \N__16180\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__16189\,
            I => \N__16177\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__16186\,
            I => \N__16174\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__16183\,
            I => \N__16171\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16167\
        );

    \I__2860\ : CascadeBuf
    port map (
            O => \N__16177\,
            I => \N__16164\
        );

    \I__2859\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16161\
        );

    \I__2858\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16158\
        );

    \I__2857\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16155\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16152\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__16164\,
            I => \N__16149\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__16161\,
            I => \N__16146\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__16158\,
            I => \N__16143\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__16155\,
            I => \N__16138\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__16152\,
            I => \N__16138\
        );

    \I__2850\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16135\
        );

    \I__2849\ : Span4Mux_s2_v
    port map (
            O => \N__16146\,
            I => \N__16132\
        );

    \I__2848\ : Span4Mux_s1_v
    port map (
            O => \N__16143\,
            I => \N__16125\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__16138\,
            I => \N__16125\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16125\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__16132\,
            I => \N__16122\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__16122\,
            I => \N__16116\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__16119\,
            I => \N__16113\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__16116\,
            I => addr_out_7
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__16113\,
            I => addr_out_7
        );

    \I__2839\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16105\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__16105\,
            I => \N__16100\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__16104\,
            I => \N__16096\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__16103\,
            I => \N__16093\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__16100\,
            I => \N__16090\
        );

    \I__2834\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16083\
        );

    \I__2833\ : InMux
    port map (
            O => \N__16096\,
            I => \N__16083\
        );

    \I__2832\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16083\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__16090\,
            I => \sb_translator_1.cnt_RNILAHE_2Z0Z_10\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__16083\,
            I => \sb_translator_1.cnt_RNILAHE_2Z0Z_10\
        );

    \I__2829\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16072\
        );

    \I__2828\ : InMux
    port map (
            O => \N__16077\,
            I => \N__16072\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16067\
        );

    \I__2826\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16062\
        );

    \I__2825\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16062\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__16067\,
            I => \N__16057\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__16062\,
            I => \N__16057\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__16057\,
            I => \sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16050\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__16053\,
            I => \N__16046\
        );

    \I__2819\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16039\
        );

    \I__2818\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16039\
        );

    \I__2817\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16039\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__16039\,
            I => \N__16035\
        );

    \I__2815\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16032\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__16035\,
            I => \N__16027\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__16032\,
            I => \N__16027\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__16027\,
            I => \sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10\
        );

    \I__2811\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16019\
        );

    \I__2810\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16016\
        );

    \I__2809\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16013\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__16019\,
            I => \N__16010\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__16016\,
            I => mosi_data_out_0
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__16013\,
            I => mosi_data_out_0
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__16010\,
            I => mosi_data_out_0
        );

    \I__2804\ : InMux
    port map (
            O => \N__16003\,
            I => \N__16000\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__16000\,
            I => \sb_translator_1.instr_tmpZ1Z_0\
        );

    \I__2802\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15993\
        );

    \I__2801\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15990\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15986\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15983\
        );

    \I__2798\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15980\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__15986\,
            I => \N__15973\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__15983\,
            I => \N__15973\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15980\,
            I => \N__15973\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__15970\,
            I => mosi_data_out_1
        );

    \I__2792\ : InMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__15964\,
            I => \sb_translator_1.instr_tmpZ1Z_1\
        );

    \I__2790\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15958\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__15958\,
            I => \N__15953\
        );

    \I__2788\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15950\
        );

    \I__2787\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15947\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__15953\,
            I => mosi_data_out_2
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__15950\,
            I => mosi_data_out_2
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__15947\,
            I => mosi_data_out_2
        );

    \I__2783\ : InMux
    port map (
            O => \N__15940\,
            I => \N__15937\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__15937\,
            I => \sb_translator_1.instr_tmpZ1Z_2\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__15934\,
            I => \N__15929\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__15933\,
            I => \N__15925\
        );

    \I__2779\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15918\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15918\
        );

    \I__2777\ : InMux
    port map (
            O => \N__15928\,
            I => \N__15913\
        );

    \I__2776\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15913\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15908\
        );

    \I__2774\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15908\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__15918\,
            I => \sb_translator_1.num_ledsZ0Z_9\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__15913\,
            I => \sb_translator_1.num_ledsZ0Z_9\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15908\,
            I => \sb_translator_1.num_ledsZ0Z_9\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \N__15897\
        );

    \I__2769\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15888\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15888\
        );

    \I__2767\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15879\
        );

    \I__2766\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15879\
        );

    \I__2765\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15879\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15879\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__15888\,
            I => \sb_translator_1.num_ledsZ0Z_11\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__15879\,
            I => \sb_translator_1.num_ledsZ0Z_11\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__15874\,
            I => \N__15869\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__15873\,
            I => \N__15864\
        );

    \I__2759\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15858\
        );

    \I__2758\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15858\
        );

    \I__2757\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15849\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15849\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15849\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15849\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__15858\,
            I => \sb_translator_1.num_ledsZ0Z_10\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__15849\,
            I => \sb_translator_1.num_ledsZ0Z_10\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__15844\,
            I => \sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_\
        );

    \I__2750\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15837\
        );

    \I__2749\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15834\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__15837\,
            I => \N__15831\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__15831\,
            I => \N__15823\
        );

    \I__2745\ : Span4Mux_v
    port map (
            O => \N__15828\,
            I => \N__15823\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__15823\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_0_0_7\
        );

    \I__2743\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15815\
        );

    \I__2742\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15810\
        );

    \I__2741\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15810\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__15815\,
            I => \N__15804\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__15810\,
            I => \N__15804\
        );

    \I__2738\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15801\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__15804\,
            I => \N__15796\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__15801\,
            I => \N__15796\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__15796\,
            I => \N__15793\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__15793\,
            I => \sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10\
        );

    \I__2733\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15787\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__15787\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_0\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__15784\,
            I => \N__15781\
        );

    \I__2730\ : CascadeBuf
    port map (
            O => \N__15781\,
            I => \N__15777\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__15780\,
            I => \N__15774\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__15777\,
            I => \N__15770\
        );

    \I__2727\ : CascadeBuf
    port map (
            O => \N__15774\,
            I => \N__15767\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__15773\,
            I => \N__15763\
        );

    \I__2725\ : CascadeBuf
    port map (
            O => \N__15770\,
            I => \N__15760\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__15767\,
            I => \N__15757\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__15766\,
            I => \N__15754\
        );

    \I__2722\ : CascadeBuf
    port map (
            O => \N__15763\,
            I => \N__15751\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__15760\,
            I => \N__15748\
        );

    \I__2720\ : CascadeBuf
    port map (
            O => \N__15757\,
            I => \N__15745\
        );

    \I__2719\ : CascadeBuf
    port map (
            O => \N__15754\,
            I => \N__15742\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__15751\,
            I => \N__15739\
        );

    \I__2717\ : CascadeBuf
    port map (
            O => \N__15748\,
            I => \N__15736\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__15745\,
            I => \N__15733\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__15742\,
            I => \N__15730\
        );

    \I__2714\ : CascadeBuf
    port map (
            O => \N__15739\,
            I => \N__15727\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__15736\,
            I => \N__15724\
        );

    \I__2712\ : CascadeBuf
    port map (
            O => \N__15733\,
            I => \N__15721\
        );

    \I__2711\ : CascadeBuf
    port map (
            O => \N__15730\,
            I => \N__15718\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__15727\,
            I => \N__15715\
        );

    \I__2709\ : CascadeBuf
    port map (
            O => \N__15724\,
            I => \N__15712\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__15721\,
            I => \N__15709\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__15718\,
            I => \N__15706\
        );

    \I__2706\ : CascadeBuf
    port map (
            O => \N__15715\,
            I => \N__15703\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__15712\,
            I => \N__15700\
        );

    \I__2704\ : CascadeBuf
    port map (
            O => \N__15709\,
            I => \N__15697\
        );

    \I__2703\ : CascadeBuf
    port map (
            O => \N__15706\,
            I => \N__15694\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__15703\,
            I => \N__15691\
        );

    \I__2701\ : CascadeBuf
    port map (
            O => \N__15700\,
            I => \N__15688\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__15697\,
            I => \N__15685\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__15694\,
            I => \N__15682\
        );

    \I__2698\ : CascadeBuf
    port map (
            O => \N__15691\,
            I => \N__15679\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__15688\,
            I => \N__15676\
        );

    \I__2696\ : CascadeBuf
    port map (
            O => \N__15685\,
            I => \N__15673\
        );

    \I__2695\ : CascadeBuf
    port map (
            O => \N__15682\,
            I => \N__15670\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \N__15667\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__15676\,
            I => \N__15664\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__15673\,
            I => \N__15661\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \N__15658\
        );

    \I__2690\ : CascadeBuf
    port map (
            O => \N__15667\,
            I => \N__15655\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__15664\,
            I => \N__15652\
        );

    \I__2688\ : CascadeBuf
    port map (
            O => \N__15661\,
            I => \N__15649\
        );

    \I__2687\ : CascadeBuf
    port map (
            O => \N__15658\,
            I => \N__15646\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__15655\,
            I => \N__15643\
        );

    \I__2685\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15640\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15637\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \N__15634\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__15643\,
            I => \N__15631\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__15640\,
            I => \N__15628\
        );

    \I__2680\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15625\
        );

    \I__2679\ : CascadeBuf
    port map (
            O => \N__15634\,
            I => \N__15622\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__15631\,
            I => \N__15618\
        );

    \I__2677\ : Span4Mux_s1_v
    port map (
            O => \N__15628\,
            I => \N__15615\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15612\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__15622\,
            I => \N__15609\
        );

    \I__2674\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15606\
        );

    \I__2673\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15603\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__15615\,
            I => \N__15598\
        );

    \I__2671\ : Span4Mux_s1_v
    port map (
            O => \N__15612\,
            I => \N__15598\
        );

    \I__2670\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15595\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__15606\,
            I => \N__15592\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__15603\,
            I => \N__15589\
        );

    \I__2667\ : Sp12to4
    port map (
            O => \N__15598\,
            I => \N__15584\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15584\
        );

    \I__2665\ : Span12Mux_s9_v
    port map (
            O => \N__15592\,
            I => \N__15581\
        );

    \I__2664\ : Span12Mux_s7_h
    port map (
            O => \N__15589\,
            I => \N__15576\
        );

    \I__2663\ : Span12Mux_s6_h
    port map (
            O => \N__15584\,
            I => \N__15576\
        );

    \I__2662\ : Odrv12
    port map (
            O => \N__15581\,
            I => addr_out_0
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__15576\,
            I => addr_out_0
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__15571\,
            I => \N__15568\
        );

    \I__2659\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15565\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__15565\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_1\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__15562\,
            I => \N__15558\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__15561\,
            I => \N__15555\
        );

    \I__2655\ : CascadeBuf
    port map (
            O => \N__15558\,
            I => \N__15550\
        );

    \I__2654\ : CascadeBuf
    port map (
            O => \N__15555\,
            I => \N__15547\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__15554\,
            I => \N__15544\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__15553\,
            I => \N__15541\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__15550\,
            I => \N__15538\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__15547\,
            I => \N__15535\
        );

    \I__2649\ : CascadeBuf
    port map (
            O => \N__15544\,
            I => \N__15532\
        );

    \I__2648\ : CascadeBuf
    port map (
            O => \N__15541\,
            I => \N__15529\
        );

    \I__2647\ : CascadeBuf
    port map (
            O => \N__15538\,
            I => \N__15526\
        );

    \I__2646\ : CascadeBuf
    port map (
            O => \N__15535\,
            I => \N__15523\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__15532\,
            I => \N__15520\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15517\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__15526\,
            I => \N__15514\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__15523\,
            I => \N__15511\
        );

    \I__2641\ : CascadeBuf
    port map (
            O => \N__15520\,
            I => \N__15508\
        );

    \I__2640\ : CascadeBuf
    port map (
            O => \N__15517\,
            I => \N__15505\
        );

    \I__2639\ : CascadeBuf
    port map (
            O => \N__15514\,
            I => \N__15502\
        );

    \I__2638\ : CascadeBuf
    port map (
            O => \N__15511\,
            I => \N__15499\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__15508\,
            I => \N__15496\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__15505\,
            I => \N__15493\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__15502\,
            I => \N__15490\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__15499\,
            I => \N__15487\
        );

    \I__2633\ : CascadeBuf
    port map (
            O => \N__15496\,
            I => \N__15484\
        );

    \I__2632\ : CascadeBuf
    port map (
            O => \N__15493\,
            I => \N__15481\
        );

    \I__2631\ : CascadeBuf
    port map (
            O => \N__15490\,
            I => \N__15478\
        );

    \I__2630\ : CascadeBuf
    port map (
            O => \N__15487\,
            I => \N__15475\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__15484\,
            I => \N__15472\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__15481\,
            I => \N__15469\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__15478\,
            I => \N__15466\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__15475\,
            I => \N__15463\
        );

    \I__2625\ : CascadeBuf
    port map (
            O => \N__15472\,
            I => \N__15460\
        );

    \I__2624\ : CascadeBuf
    port map (
            O => \N__15469\,
            I => \N__15457\
        );

    \I__2623\ : CascadeBuf
    port map (
            O => \N__15466\,
            I => \N__15454\
        );

    \I__2622\ : CascadeBuf
    port map (
            O => \N__15463\,
            I => \N__15451\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__15460\,
            I => \N__15448\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__15457\,
            I => \N__15445\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__15454\,
            I => \N__15442\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15439\
        );

    \I__2617\ : CascadeBuf
    port map (
            O => \N__15448\,
            I => \N__15436\
        );

    \I__2616\ : CascadeBuf
    port map (
            O => \N__15445\,
            I => \N__15433\
        );

    \I__2615\ : CascadeBuf
    port map (
            O => \N__15442\,
            I => \N__15430\
        );

    \I__2614\ : CascadeBuf
    port map (
            O => \N__15439\,
            I => \N__15427\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__15436\,
            I => \N__15424\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__15433\,
            I => \N__15421\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__15430\,
            I => \N__15418\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__15427\,
            I => \N__15415\
        );

    \I__2609\ : CascadeBuf
    port map (
            O => \N__15424\,
            I => \N__15412\
        );

    \I__2608\ : CascadeBuf
    port map (
            O => \N__15421\,
            I => \N__15409\
        );

    \I__2607\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15405\
        );

    \I__2606\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15402\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \N__15399\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15396\
        );

    \I__2603\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15393\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__15405\,
            I => \N__15388\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__15402\,
            I => \N__15388\
        );

    \I__2600\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15385\
        );

    \I__2599\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15382\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__15393\,
            I => \N__15379\
        );

    \I__2597\ : Span4Mux_s3_v
    port map (
            O => \N__15388\,
            I => \N__15376\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15371\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15371\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__15379\,
            I => \N__15364\
        );

    \I__2593\ : Span4Mux_h
    port map (
            O => \N__15376\,
            I => \N__15364\
        );

    \I__2592\ : Span4Mux_s3_v
    port map (
            O => \N__15371\,
            I => \N__15364\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__15364\,
            I => \N__15361\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__15361\,
            I => \N__15358\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__15358\,
            I => addr_out_1
        );

    \I__2588\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15352\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__15352\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_2\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__15349\,
            I => \N__15346\
        );

    \I__2585\ : CascadeBuf
    port map (
            O => \N__15346\,
            I => \N__15343\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__15343\,
            I => \N__15338\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__15342\,
            I => \N__15335\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \N__15332\
        );

    \I__2581\ : CascadeBuf
    port map (
            O => \N__15338\,
            I => \N__15329\
        );

    \I__2580\ : CascadeBuf
    port map (
            O => \N__15335\,
            I => \N__15326\
        );

    \I__2579\ : CascadeBuf
    port map (
            O => \N__15332\,
            I => \N__15322\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__15329\,
            I => \N__15319\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__15326\,
            I => \N__15316\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15313\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__15322\,
            I => \N__15310\
        );

    \I__2574\ : CascadeBuf
    port map (
            O => \N__15319\,
            I => \N__15307\
        );

    \I__2573\ : CascadeBuf
    port map (
            O => \N__15316\,
            I => \N__15304\
        );

    \I__2572\ : CascadeBuf
    port map (
            O => \N__15313\,
            I => \N__15301\
        );

    \I__2571\ : CascadeBuf
    port map (
            O => \N__15310\,
            I => \N__15298\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__15307\,
            I => \N__15295\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__15304\,
            I => \N__15292\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__15301\,
            I => \N__15289\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__15298\,
            I => \N__15286\
        );

    \I__2566\ : CascadeBuf
    port map (
            O => \N__15295\,
            I => \N__15283\
        );

    \I__2565\ : CascadeBuf
    port map (
            O => \N__15292\,
            I => \N__15280\
        );

    \I__2564\ : CascadeBuf
    port map (
            O => \N__15289\,
            I => \N__15277\
        );

    \I__2563\ : CascadeBuf
    port map (
            O => \N__15286\,
            I => \N__15274\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__15283\,
            I => \N__15271\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \N__15268\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__15277\,
            I => \N__15265\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \N__15262\
        );

    \I__2558\ : CascadeBuf
    port map (
            O => \N__15271\,
            I => \N__15259\
        );

    \I__2557\ : CascadeBuf
    port map (
            O => \N__15268\,
            I => \N__15256\
        );

    \I__2556\ : CascadeBuf
    port map (
            O => \N__15265\,
            I => \N__15253\
        );

    \I__2555\ : CascadeBuf
    port map (
            O => \N__15262\,
            I => \N__15250\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__15259\,
            I => \N__15247\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__15256\,
            I => \N__15244\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__15253\,
            I => \N__15241\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__15250\,
            I => \N__15238\
        );

    \I__2550\ : CascadeBuf
    port map (
            O => \N__15247\,
            I => \N__15235\
        );

    \I__2549\ : CascadeBuf
    port map (
            O => \N__15244\,
            I => \N__15232\
        );

    \I__2548\ : CascadeBuf
    port map (
            O => \N__15241\,
            I => \N__15229\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__15238\,
            I => \N__15226\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__15235\,
            I => \N__15223\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__15232\,
            I => \N__15220\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__15229\,
            I => \N__15217\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__15226\,
            I => \N__15214\
        );

    \I__2542\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15211\
        );

    \I__2541\ : CascadeBuf
    port map (
            O => \N__15220\,
            I => \N__15208\
        );

    \I__2540\ : CascadeBuf
    port map (
            O => \N__15217\,
            I => \N__15205\
        );

    \I__2539\ : CascadeBuf
    port map (
            O => \N__15214\,
            I => \N__15202\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15199\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__15208\,
            I => \N__15196\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \N__15193\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__15202\,
            I => \N__15190\
        );

    \I__2534\ : Span4Mux_s1_v
    port map (
            O => \N__15199\,
            I => \N__15186\
        );

    \I__2533\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15183\
        );

    \I__2532\ : CascadeBuf
    port map (
            O => \N__15193\,
            I => \N__15180\
        );

    \I__2531\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15177\
        );

    \I__2530\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15174\
        );

    \I__2529\ : Span4Mux_s2_h
    port map (
            O => \N__15186\,
            I => \N__15169\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__15183\,
            I => \N__15169\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__15180\,
            I => \N__15166\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15163\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15158\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__15169\,
            I => \N__15158\
        );

    \I__2523\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15155\
        );

    \I__2522\ : Span4Mux_s1_v
    port map (
            O => \N__15163\,
            I => \N__15148\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__15158\,
            I => \N__15148\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__15155\,
            I => \N__15148\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__15148\,
            I => \N__15145\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__15145\,
            I => \N__15142\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__15142\,
            I => addr_out_2
        );

    \I__2516\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15136\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__15136\,
            I => \N__15133\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__15133\,
            I => \sb_translator_1.addr_out_RNO_0Z0Z_3\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__15130\,
            I => \N__15125\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__15129\,
            I => \N__15121\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__15128\,
            I => \N__15118\
        );

    \I__2510\ : CascadeBuf
    port map (
            O => \N__15125\,
            I => \N__15115\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__15124\,
            I => \N__15112\
        );

    \I__2508\ : CascadeBuf
    port map (
            O => \N__15121\,
            I => \N__15109\
        );

    \I__2507\ : CascadeBuf
    port map (
            O => \N__15118\,
            I => \N__15106\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__15115\,
            I => \N__15103\
        );

    \I__2505\ : CascadeBuf
    port map (
            O => \N__15112\,
            I => \N__15100\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__15109\,
            I => \N__15097\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__15106\,
            I => \N__15094\
        );

    \I__2502\ : CascadeBuf
    port map (
            O => \N__15103\,
            I => \N__15091\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__15100\,
            I => \N__15088\
        );

    \I__2500\ : CascadeBuf
    port map (
            O => \N__15097\,
            I => \N__15085\
        );

    \I__2499\ : CascadeBuf
    port map (
            O => \N__15094\,
            I => \N__15082\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__15091\,
            I => \N__15079\
        );

    \I__2497\ : CascadeBuf
    port map (
            O => \N__15088\,
            I => \N__15076\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__15085\,
            I => \N__15073\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \N__15070\
        );

    \I__2494\ : CascadeBuf
    port map (
            O => \N__15079\,
            I => \N__15067\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__15076\,
            I => \N__15064\
        );

    \I__2492\ : CascadeBuf
    port map (
            O => \N__15073\,
            I => \N__15061\
        );

    \I__2491\ : CascadeBuf
    port map (
            O => \N__15070\,
            I => \N__15058\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__15067\,
            I => \N__15055\
        );

    \I__2489\ : CascadeBuf
    port map (
            O => \N__15064\,
            I => \N__15052\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__15061\,
            I => \N__15049\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__15058\,
            I => \N__15046\
        );

    \I__2486\ : CascadeBuf
    port map (
            O => \N__15055\,
            I => \N__15043\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__15052\,
            I => \N__15040\
        );

    \I__2484\ : CascadeBuf
    port map (
            O => \N__15049\,
            I => \N__15037\
        );

    \I__2483\ : CascadeBuf
    port map (
            O => \N__15046\,
            I => \N__15034\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__15043\,
            I => \N__15031\
        );

    \I__2481\ : CascadeBuf
    port map (
            O => \N__15040\,
            I => \N__15028\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__15037\,
            I => \N__15025\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__15034\,
            I => \N__15022\
        );

    \I__2478\ : CascadeBuf
    port map (
            O => \N__15031\,
            I => \N__15019\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__15028\,
            I => \N__15016\
        );

    \I__2476\ : CascadeBuf
    port map (
            O => \N__15025\,
            I => \N__15013\
        );

    \I__2475\ : CascadeBuf
    port map (
            O => \N__15022\,
            I => \N__15010\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__15019\,
            I => \N__15007\
        );

    \I__2473\ : CascadeBuf
    port map (
            O => \N__15016\,
            I => \N__15004\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \N__15001\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__15010\,
            I => \N__14998\
        );

    \I__2470\ : CascadeBuf
    port map (
            O => \N__15007\,
            I => \N__14995\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__15004\,
            I => \N__14992\
        );

    \I__2468\ : CascadeBuf
    port map (
            O => \N__15001\,
            I => \N__14989\
        );

    \I__2467\ : CascadeBuf
    port map (
            O => \N__14998\,
            I => \N__14986\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__14995\,
            I => \N__14983\
        );

    \I__2465\ : CascadeBuf
    port map (
            O => \N__14992\,
            I => \N__14980\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \N__14977\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__14986\,
            I => \N__14974\
        );

    \I__2462\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14970\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__14980\,
            I => \N__14967\
        );

    \I__2460\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14964\
        );

    \I__2459\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14961\
        );

    \I__2458\ : InMux
    port map (
            O => \N__14973\,
            I => \N__14958\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__14970\,
            I => \N__14955\
        );

    \I__2456\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14952\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__14964\,
            I => \N__14949\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__14961\,
            I => \N__14946\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__14958\,
            I => \N__14941\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__14955\,
            I => \N__14941\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__14952\,
            I => \N__14938\
        );

    \I__2450\ : Span4Mux_h
    port map (
            O => \N__14949\,
            I => \N__14933\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__14946\,
            I => \N__14933\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__14941\,
            I => \N__14928\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__14938\,
            I => \N__14928\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__14933\,
            I => \N__14925\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__14928\,
            I => \N__14922\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__14925\,
            I => \N__14919\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__14922\,
            I => \N__14916\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__14919\,
            I => addr_out_3
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__14916\,
            I => addr_out_3
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__14911\,
            I => \N__14908\
        );

    \I__2439\ : CascadeBuf
    port map (
            O => \N__14908\,
            I => \N__14902\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__14907\,
            I => \N__14899\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__14906\,
            I => \N__14896\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \N__14893\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__14902\,
            I => \N__14890\
        );

    \I__2434\ : CascadeBuf
    port map (
            O => \N__14899\,
            I => \N__14887\
        );

    \I__2433\ : CascadeBuf
    port map (
            O => \N__14896\,
            I => \N__14884\
        );

    \I__2432\ : CascadeBuf
    port map (
            O => \N__14893\,
            I => \N__14881\
        );

    \I__2431\ : CascadeBuf
    port map (
            O => \N__14890\,
            I => \N__14878\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__14887\,
            I => \N__14875\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__14884\,
            I => \N__14872\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__14881\,
            I => \N__14869\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__14878\,
            I => \N__14866\
        );

    \I__2426\ : CascadeBuf
    port map (
            O => \N__14875\,
            I => \N__14863\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__14872\,
            I => \N__14860\
        );

    \I__2424\ : CascadeBuf
    port map (
            O => \N__14869\,
            I => \N__14857\
        );

    \I__2423\ : CascadeBuf
    port map (
            O => \N__14866\,
            I => \N__14854\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__14863\,
            I => \N__14851\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__14860\,
            I => \N__14848\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__14857\,
            I => \N__14845\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__14854\,
            I => \N__14842\
        );

    \I__2418\ : CascadeBuf
    port map (
            O => \N__14851\,
            I => \N__14839\
        );

    \I__2417\ : CascadeBuf
    port map (
            O => \N__14848\,
            I => \N__14836\
        );

    \I__2416\ : CascadeBuf
    port map (
            O => \N__14845\,
            I => \N__14833\
        );

    \I__2415\ : CascadeBuf
    port map (
            O => \N__14842\,
            I => \N__14830\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__14839\,
            I => \N__14827\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__14836\,
            I => \N__14824\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__14833\,
            I => \N__14821\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__14830\,
            I => \N__14818\
        );

    \I__2410\ : CascadeBuf
    port map (
            O => \N__14827\,
            I => \N__14815\
        );

    \I__2409\ : CascadeBuf
    port map (
            O => \N__14824\,
            I => \N__14812\
        );

    \I__2408\ : CascadeBuf
    port map (
            O => \N__14821\,
            I => \N__14809\
        );

    \I__2407\ : CascadeBuf
    port map (
            O => \N__14818\,
            I => \N__14806\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14803\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__14812\,
            I => \N__14800\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__14809\,
            I => \N__14797\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__14806\,
            I => \N__14794\
        );

    \I__2402\ : CascadeBuf
    port map (
            O => \N__14803\,
            I => \N__14791\
        );

    \I__2401\ : CascadeBuf
    port map (
            O => \N__14800\,
            I => \N__14788\
        );

    \I__2400\ : CascadeBuf
    port map (
            O => \N__14797\,
            I => \N__14785\
        );

    \I__2399\ : CascadeBuf
    port map (
            O => \N__14794\,
            I => \N__14782\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__14791\,
            I => \N__14779\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__14788\,
            I => \N__14776\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__14785\,
            I => \N__14773\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__14782\,
            I => \N__14770\
        );

    \I__2394\ : CascadeBuf
    port map (
            O => \N__14779\,
            I => \N__14766\
        );

    \I__2393\ : CascadeBuf
    port map (
            O => \N__14776\,
            I => \N__14763\
        );

    \I__2392\ : CascadeBuf
    port map (
            O => \N__14773\,
            I => \N__14760\
        );

    \I__2391\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14757\
        );

    \I__2390\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14754\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__14766\,
            I => \N__14751\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__14763\,
            I => \N__14748\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__14760\,
            I => \N__14745\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__14757\,
            I => \N__14742\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__14754\,
            I => \N__14739\
        );

    \I__2384\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14736\
        );

    \I__2383\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14733\
        );

    \I__2382\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14730\
        );

    \I__2381\ : Span4Mux_s1_v
    port map (
            O => \N__14742\,
            I => \N__14727\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__14739\,
            I => \N__14722\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__14736\,
            I => \N__14722\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__14733\,
            I => \N__14717\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__14730\,
            I => \N__14717\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__14727\,
            I => \N__14712\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__14722\,
            I => \N__14712\
        );

    \I__2374\ : Span12Mux_s9_v
    port map (
            O => \N__14717\,
            I => \N__14709\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__14712\,
            I => \N__14706\
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__14709\,
            I => addr_out_4
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__14706\,
            I => addr_out_4
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__14701\,
            I => \sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_\
        );

    \I__2369\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__14695\,
            I => miso_data_in_13
        );

    \I__2367\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14689\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__14689\,
            I => miso_data_in_14
        );

    \I__2365\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14683\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__14683\,
            I => miso_data_in_15
        );

    \I__2363\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14677\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__14677\,
            I => miso_data_in_16
        );

    \I__2361\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14668\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__14668\,
            I => \N__14664\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__14667\,
            I => \N__14661\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__14664\,
            I => \N__14658\
        );

    \I__2356\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14655\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__14658\,
            I => \sb_translator_1.instr_tmpZ0Z_17\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__14655\,
            I => \sb_translator_1.instr_tmpZ0Z_17\
        );

    \I__2353\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__14647\,
            I => miso_data_in_17
        );

    \I__2351\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14640\
        );

    \I__2350\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14637\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__14640\,
            I => mosi_data_out_11
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__14637\,
            I => mosi_data_out_11
        );

    \I__2347\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__14629\,
            I => \N__14625\
        );

    \I__2345\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14621\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__14625\,
            I => \N__14618\
        );

    \I__2343\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14615\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__14621\,
            I => \N__14612\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__14618\,
            I => \sb_translator_1.cntZ0Z_3\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__14615\,
            I => \sb_translator_1.cntZ0Z_3\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__14612\,
            I => \sb_translator_1.cntZ0Z_3\
        );

    \I__2338\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14601\
        );

    \I__2337\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14598\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__14601\,
            I => mosi_data_out_13
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__14598\,
            I => mosi_data_out_13
        );

    \I__2334\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14590\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__14590\,
            I => \N__14586\
        );

    \I__2332\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14582\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__14586\,
            I => \N__14579\
        );

    \I__2330\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14576\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__14582\,
            I => \N__14573\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__14579\,
            I => \sb_translator_1.cntZ0Z_5\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__14576\,
            I => \sb_translator_1.cntZ0Z_5\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__14573\,
            I => \sb_translator_1.cntZ0Z_5\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__2324\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__14554\,
            I => \spi_slave_1.miso_data_outZ0Z_17\
        );

    \I__2320\ : CEMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__14548\,
            I => \N__14543\
        );

    \I__2318\ : CEMux
    port map (
            O => \N__14547\,
            I => \N__14540\
        );

    \I__2317\ : CEMux
    port map (
            O => \N__14546\,
            I => \N__14536\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__14543\,
            I => \N__14531\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14531\
        );

    \I__2314\ : CEMux
    port map (
            O => \N__14539\,
            I => \N__14528\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14525\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__14531\,
            I => \N__14520\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__14528\,
            I => \N__14520\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__14525\,
            I => \N__14517\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__14520\,
            I => \N__14514\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__14517\,
            I => \spi_slave_1.bitcnt_tx_0_sqmuxa\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__14514\,
            I => \spi_slave_1.bitcnt_tx_0_sqmuxa\
        );

    \I__2306\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14506\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__14506\,
            I => miso_data_in_10
        );

    \I__2304\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14500\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__14500\,
            I => miso_data_in_11
        );

    \I__2302\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14494\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__14494\,
            I => miso_data_in_12
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__14491\,
            I => \demux.N_236_cascade_\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__14488\,
            I => \demux.N_235_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__2297\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14479\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__2295\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14463\
        );

    \I__2294\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14463\
        );

    \I__2293\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14463\
        );

    \I__2292\ : Span4Mux_h
    port map (
            O => \N__14473\,
            I => \N__14460\
        );

    \I__2291\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14453\
        );

    \I__2290\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14453\
        );

    \I__2289\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14453\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__14463\,
            I => \N__14450\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__14460\,
            I => \demux.N_424_i_0_a2Z0Z_6\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__14453\,
            I => \demux.N_424_i_0_a2Z0Z_6\
        );

    \I__2285\ : Odrv12
    port map (
            O => \N__14450\,
            I => \demux.N_424_i_0_a2Z0Z_6\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14439\
        );

    \I__2283\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14425\
        );

    \I__2282\ : InMux
    port map (
            O => \N__14439\,
            I => \N__14425\
        );

    \I__2281\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14425\
        );

    \I__2280\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14425\
        );

    \I__2279\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14425\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__14425\,
            I => \N__14422\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__14422\,
            I => ram_sel_6
        );

    \I__2276\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14404\
        );

    \I__2275\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14404\
        );

    \I__2274\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14404\
        );

    \I__2273\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14404\
        );

    \I__2272\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14404\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__14401\,
            I => ram_sel_9
        );

    \I__2269\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14395\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__2267\ : Span4Mux_s3_v
    port map (
            O => \N__14392\,
            I => \N__14389\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__14389\,
            I => \N__14386\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__14386\,
            I => miso_data_in_9
        );

    \I__2264\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14380\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__14380\,
            I => \N__14377\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__14377\,
            I => \N__14374\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__14374\,
            I => demux_data_in_56
        );

    \I__2260\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14368\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__14368\,
            I => \demux.N_424_i_0_a3Z0Z_1\
        );

    \I__2258\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14356\
        );

    \I__2257\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14356\
        );

    \I__2256\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14356\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14353\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__14353\,
            I => \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__2252\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14338\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14333\
        );

    \I__2250\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14333\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14324\
        );

    \I__2248\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14324\
        );

    \I__2247\ : InMux
    port map (
            O => \N__14342\,
            I => \N__14324\
        );

    \I__2246\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14324\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__14338\,
            I => \N__14319\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__14333\,
            I => \N__14319\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__14324\,
            I => \sb_translator_1.state_RNIHS98Z0Z_0\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__14319\,
            I => \sb_translator_1.state_RNIHS98Z0Z_0\
        );

    \I__2241\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14299\
        );

    \I__2240\ : InMux
    port map (
            O => \N__14313\,
            I => \N__14299\
        );

    \I__2239\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14299\
        );

    \I__2238\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14299\
        );

    \I__2237\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14299\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__14299\,
            I => \N__14296\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__14296\,
            I => \N__14292\
        );

    \I__2234\ : InMux
    port map (
            O => \N__14295\,
            I => \N__14289\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__14292\,
            I => \sb_translator_1.state_RNIHS98_0Z0Z_0\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__14289\,
            I => \sb_translator_1.state_RNIHS98_0Z0Z_0\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__2230\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14275\
        );

    \I__2229\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14272\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__14281\,
            I => \N__14269\
        );

    \I__2227\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14266\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14261\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14261\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14258\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14255\
        );

    \I__2222\ : Span4Mux_h
    port map (
            O => \N__14261\,
            I => \N__14252\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__14258\,
            I => \N__14249\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__14255\,
            I => \N__14246\
        );

    \I__2219\ : Span4Mux_s2_h
    port map (
            O => \N__14252\,
            I => \N__14243\
        );

    \I__2218\ : Span4Mux_h
    port map (
            O => \N__14249\,
            I => \N__14240\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__14246\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__14243\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__14240\,
            I => \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14229\
        );

    \I__2213\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14224\
        );

    \I__2212\ : InMux
    port map (
            O => \N__14229\,
            I => \N__14224\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14221\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__14221\,
            I => \sb_translator_1.N_1089\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14212\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__14212\,
            I => \N__14209\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__14209\,
            I => \N__14206\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__14206\,
            I => \N__14203\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__14203\,
            I => demux_data_in_74
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__14200\,
            I => \N__14197\
        );

    \I__2202\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14194\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__14194\,
            I => \N__14191\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__14191\,
            I => \N__14188\
        );

    \I__2199\ : Span4Mux_h
    port map (
            O => \N__14188\,
            I => \N__14185\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__14185\,
            I => demux_data_in_82
        );

    \I__2197\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14179\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N__14176\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__14176\,
            I => \N__14173\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__14173\,
            I => demux_data_in_50
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__14170\,
            I => \demux.N_422_i_0_o2Z0Z_6_cascade_\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14164\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__14164\,
            I => \N__14161\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__14161\,
            I => \N__14158\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__14155\,
            I => demux_data_in_73
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__14152\,
            I => \N__14149\
        );

    \I__2186\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14146\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__14146\,
            I => \N__14143\
        );

    \I__2184\ : Span12Mux_s10_h
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__2183\ : Odrv12
    port map (
            O => \N__14140\,
            I => demux_data_in_81
        );

    \I__2182\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14134\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__14134\,
            I => \N__14131\
        );

    \I__2180\ : Span4Mux_v
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__14128\,
            I => demux_data_in_49
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__14125\,
            I => \demux.N_423_i_0_o2Z0Z_6_cascade_\
        );

    \I__2177\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14119\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__14119\,
            I => \demux.N_423_i_0_a3Z0Z_1\
        );

    \I__2175\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14113\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__14113\,
            I => \N__14110\
        );

    \I__2173\ : Span4Mux_h
    port map (
            O => \N__14110\,
            I => \N__14107\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__14107\,
            I => demux_data_in_58
        );

    \I__2171\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14101\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__14101\,
            I => \demux.N_422_i_0_a3Z0Z_1\
        );

    \I__2169\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__14095\,
            I => \N__14092\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__14092\,
            I => \N__14089\
        );

    \I__2166\ : Span4Mux_h
    port map (
            O => \N__14089\,
            I => \N__14086\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__14086\,
            I => demux_data_in_80
        );

    \I__2164\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14080\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__14080\,
            I => \N__14077\
        );

    \I__2162\ : Span12Mux_s10_h
    port map (
            O => \N__14077\,
            I => \N__14074\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__14074\,
            I => demux_data_in_72
        );

    \I__2160\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14068\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__14065\,
            I => \N__14062\
        );

    \I__2157\ : Span4Mux_s3_h
    port map (
            O => \N__14062\,
            I => \N__14059\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__14059\,
            I => demux_data_in_48
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__14056\,
            I => \demux.N_424_i_0_o2_6_cascade_\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__2153\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14043\
        );

    \I__2152\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__2151\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14040\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__14043\,
            I => \sb_translator_1.cnt_RNILAHE_0Z0Z_10\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__14040\,
            I => \sb_translator_1.cnt_RNILAHE_0Z0Z_10\
        );

    \I__2148\ : CEMux
    port map (
            O => \N__14035\,
            I => \N__14032\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__14026\,
            I => \N__14023\
        );

    \I__2144\ : Sp12to4
    port map (
            O => \N__14023\,
            I => \N__14020\
        );

    \I__2143\ : Span12Mux_s6_v
    port map (
            O => \N__14020\,
            I => \N__14017\
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__14017\,
            I => ram_we_4
        );

    \I__2141\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14002\
        );

    \I__2140\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14002\
        );

    \I__2139\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14002\
        );

    \I__2138\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14002\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__14002\,
            I => \N__13999\
        );

    \I__2136\ : Span4Mux_h
    port map (
            O => \N__13999\,
            I => \N__13996\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__13996\,
            I => \sb_translator_1.cnt_RNIJ7EF_2Z0Z_9\
        );

    \I__2134\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13972\
        );

    \I__2133\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13972\
        );

    \I__2132\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13972\
        );

    \I__2131\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13972\
        );

    \I__2130\ : InMux
    port map (
            O => \N__13989\,
            I => \N__13972\
        );

    \I__2129\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13972\
        );

    \I__2128\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13972\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__13972\,
            I => \sb_translator_1.state_RNI9ILJ_0Z0Z_0\
        );

    \I__2126\ : CEMux
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13963\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__13963\,
            I => \N__13960\
        );

    \I__2123\ : Sp12to4
    port map (
            O => \N__13960\,
            I => \N__13957\
        );

    \I__2122\ : Span12Mux_s7_v
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__13954\,
            I => ram_we_6
        );

    \I__2120\ : InMux
    port map (
            O => \N__13951\,
            I => \N__13948\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__2118\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13935\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13935\
        );

    \I__2116\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13935\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__13942\,
            I => \N__13932\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13935\,
            I => \N__13929\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__13932\,
            I => \sb_translator_1.cnt_RNIJ7EF_1Z0Z_9\
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__13929\,
            I => \sb_translator_1.cnt_RNIJ7EF_1Z0Z_9\
        );

    \I__2111\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13915\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13902\
        );

    \I__2109\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13902\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13902\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13902\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13902\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13902\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13915\,
            I => \sb_translator_1.state_RNI9ILJZ0Z_0\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13902\,
            I => \sb_translator_1.state_RNI9ILJZ0Z_0\
        );

    \I__2102\ : CEMux
    port map (
            O => \N__13897\,
            I => \N__13894\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2100\ : Span4Mux_s3_h
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__13882\,
            I => ram_we_1
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__13879\,
            I => \sb_translator_1.N_1091_cascade_\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__13876\,
            I => \sb_translator_1.N_1089_cascade_\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__13873\,
            I => \N__13869\
        );

    \I__2093\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13864\
        );

    \I__2092\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13864\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__13864\,
            I => \sb_translator_1.N_1091\
        );

    \I__2090\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__13858\,
            I => \sb_translator_1.instr_tmpZ1Z_5\
        );

    \I__2088\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13852\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__2086\ : Span4Mux_s1_v
    port map (
            O => \N__13849\,
            I => \N__13844\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13841\
        );

    \I__2084\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13838\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__13844\,
            I => mosi_data_out_5
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__13841\,
            I => mosi_data_out_5
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__13838\,
            I => mosi_data_out_5
        );

    \I__2080\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13827\
        );

    \I__2079\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13819\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__13827\,
            I => \N__13815\
        );

    \I__2077\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13812\
        );

    \I__2076\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13809\
        );

    \I__2075\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13806\
        );

    \I__2074\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13803\
        );

    \I__2073\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13799\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__13819\,
            I => \N__13795\
        );

    \I__2071\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13792\
        );

    \I__2070\ : Span4Mux_s3_v
    port map (
            O => \N__13815\,
            I => \N__13781\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__13812\,
            I => \N__13781\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__13809\,
            I => \N__13781\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13776\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__13803\,
            I => \N__13776\
        );

    \I__2065\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13773\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__13799\,
            I => \N__13770\
        );

    \I__2063\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13767\
        );

    \I__2062\ : Span4Mux_s3_h
    port map (
            O => \N__13795\,
            I => \N__13762\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13762\
        );

    \I__2060\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13759\
        );

    \I__2059\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13756\
        );

    \I__2058\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13753\
        );

    \I__2057\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13750\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__13781\,
            I => \N__13743\
        );

    \I__2055\ : Span4Mux_s2_v
    port map (
            O => \N__13776\,
            I => \N__13743\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__13773\,
            I => \N__13743\
        );

    \I__2053\ : Span4Mux_s0_v
    port map (
            O => \N__13770\,
            I => \N__13738\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__13767\,
            I => \N__13738\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__13762\,
            I => \N__13731\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__13759\,
            I => \N__13731\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13731\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13728\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__13750\,
            I => \N__13725\
        );

    \I__2046\ : Sp12to4
    port map (
            O => \N__13743\,
            I => \N__13722\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__13738\,
            I => \N__13713\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__13731\,
            I => \N__13713\
        );

    \I__2043\ : Span4Mux_s3_h
    port map (
            O => \N__13728\,
            I => \N__13713\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__13725\,
            I => \N__13713\
        );

    \I__2041\ : Span12Mux_s5_v
    port map (
            O => \N__13722\,
            I => \N__13710\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__13713\,
            I => \N__13707\
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__13710\,
            I => ram_data_in_5
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__13707\,
            I => ram_data_in_5
        );

    \I__2037\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13699\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__13696\,
            I => \sb_translator_1.instr_tmpZ0Z_6\
        );

    \I__2034\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__13690\,
            I => \N__13685\
        );

    \I__2032\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13682\
        );

    \I__2031\ : InMux
    port map (
            O => \N__13688\,
            I => \N__13679\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__13685\,
            I => mosi_data_out_6
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__13682\,
            I => mosi_data_out_6
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__13679\,
            I => mosi_data_out_6
        );

    \I__2027\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13666\
        );

    \I__2026\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13659\
        );

    \I__2025\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13656\
        );

    \I__2024\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13652\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__13666\,
            I => \N__13649\
        );

    \I__2022\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13646\
        );

    \I__2021\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13642\
        );

    \I__2020\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13639\
        );

    \I__2019\ : InMux
    port map (
            O => \N__13662\,
            I => \N__13635\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__13659\,
            I => \N__13631\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__13656\,
            I => \N__13628\
        );

    \I__2016\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13625\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13621\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__13649\,
            I => \N__13618\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13615\
        );

    \I__2012\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13612\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__13642\,
            I => \N__13606\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__13639\,
            I => \N__13606\
        );

    \I__2009\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13603\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13600\
        );

    \I__2007\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13597\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__13631\,
            I => \N__13594\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__13628\,
            I => \N__13591\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__13625\,
            I => \N__13588\
        );

    \I__2003\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13585\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__13621\,
            I => \N__13582\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__13618\,
            I => \N__13577\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__13615\,
            I => \N__13577\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__13612\,
            I => \N__13574\
        );

    \I__1998\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13571\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__13606\,
            I => \N__13566\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__13603\,
            I => \N__13566\
        );

    \I__1995\ : Span4Mux_s1_v
    port map (
            O => \N__13600\,
            I => \N__13561\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__13597\,
            I => \N__13561\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__13594\,
            I => \N__13554\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__13591\,
            I => \N__13554\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__13588\,
            I => \N__13554\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__13585\,
            I => \N__13551\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__13582\,
            I => \N__13544\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__13577\,
            I => \N__13544\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__13574\,
            I => \N__13544\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__13571\,
            I => \N__13541\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__13566\,
            I => \N__13536\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__13561\,
            I => \N__13536\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__13554\,
            I => \N__13531\
        );

    \I__1982\ : Span4Mux_h
    port map (
            O => \N__13551\,
            I => \N__13531\
        );

    \I__1981\ : Span4Mux_h
    port map (
            O => \N__13544\,
            I => \N__13526\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__13541\,
            I => \N__13526\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__13536\,
            I => ram_data_in_6
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__13531\,
            I => ram_data_in_6
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__13526\,
            I => ram_data_in_6
        );

    \I__1976\ : InMux
    port map (
            O => \N__13519\,
            I => \N__13516\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__13516\,
            I => \sb_translator_1.instr_tmpZ0Z_7\
        );

    \I__1974\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13505\
        );

    \I__1972\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13502\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13499\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__13505\,
            I => mosi_data_out_7
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__13502\,
            I => mosi_data_out_7
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__13499\,
            I => mosi_data_out_7
        );

    \I__1967\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13488\
        );

    \I__1966\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13481\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__13488\,
            I => \N__13478\
        );

    \I__1964\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13473\
        );

    \I__1963\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13468\
        );

    \I__1962\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13465\
        );

    \I__1961\ : InMux
    port map (
            O => \N__13484\,
            I => \N__13461\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__13481\,
            I => \N__13457\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__13478\,
            I => \N__13454\
        );

    \I__1958\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13451\
        );

    \I__1957\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13447\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__13473\,
            I => \N__13444\
        );

    \I__1955\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13441\
        );

    \I__1954\ : InMux
    port map (
            O => \N__13471\,
            I => \N__13437\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__13468\,
            I => \N__13432\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__13465\,
            I => \N__13432\
        );

    \I__1951\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13429\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__13461\,
            I => \N__13426\
        );

    \I__1949\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13423\
        );

    \I__1948\ : Span4Mux_h
    port map (
            O => \N__13457\,
            I => \N__13420\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__13454\,
            I => \N__13415\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__13451\,
            I => \N__13415\
        );

    \I__1945\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13412\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__13447\,
            I => \N__13409\
        );

    \I__1943\ : Span4Mux_h
    port map (
            O => \N__13444\,
            I => \N__13406\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__13441\,
            I => \N__13403\
        );

    \I__1941\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13400\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__13437\,
            I => \N__13397\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__13432\,
            I => \N__13392\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__13429\,
            I => \N__13392\
        );

    \I__1937\ : Span4Mux_s1_v
    port map (
            O => \N__13426\,
            I => \N__13387\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__13423\,
            I => \N__13387\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__13420\,
            I => \N__13382\
        );

    \I__1934\ : Span4Mux_h
    port map (
            O => \N__13415\,
            I => \N__13382\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__13412\,
            I => \N__13379\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__13409\,
            I => \N__13376\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__13406\,
            I => \N__13371\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__13403\,
            I => \N__13371\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__13400\,
            I => \N__13368\
        );

    \I__1928\ : Span12Mux_s8_h
    port map (
            O => \N__13397\,
            I => \N__13365\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__13392\,
            I => \N__13360\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__13387\,
            I => \N__13360\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__13382\,
            I => \N__13355\
        );

    \I__1924\ : Span4Mux_h
    port map (
            O => \N__13379\,
            I => \N__13355\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__13376\,
            I => \N__13348\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__13371\,
            I => \N__13348\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__13368\,
            I => \N__13348\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__13365\,
            I => ram_data_in_7
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__13360\,
            I => ram_data_in_7
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__13355\,
            I => ram_data_in_7
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__13348\,
            I => ram_data_in_7
        );

    \I__1916\ : CEMux
    port map (
            O => \N__13339\,
            I => \N__13336\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__13336\,
            I => \N__13333\
        );

    \I__1914\ : Span4Mux_s2_v
    port map (
            O => \N__13333\,
            I => \N__13330\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__13330\,
            I => \N__13327\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__13327\,
            I => ram_we_0
        );

    \I__1911\ : CEMux
    port map (
            O => \N__13324\,
            I => \N__13321\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13318\
        );

    \I__1909\ : Span4Mux_s1_v
    port map (
            O => \N__13318\,
            I => \N__13315\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__13315\,
            I => \N__13312\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__13312\,
            I => \N__13309\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__13309\,
            I => ram_we_2
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__13306\,
            I => \N__13303\
        );

    \I__1904\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13296\
        );

    \I__1903\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13296\
        );

    \I__1902\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13293\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__13296\,
            I => \sb_translator_1.cnt_RNILAHE_1Z0Z_10\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__13293\,
            I => \sb_translator_1.cnt_RNILAHE_1Z0Z_10\
        );

    \I__1899\ : CEMux
    port map (
            O => \N__13288\,
            I => \N__13285\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__13285\,
            I => \N__13282\
        );

    \I__1897\ : Span4Mux_s3_v
    port map (
            O => \N__13282\,
            I => \N__13279\
        );

    \I__1896\ : Span4Mux_s3_h
    port map (
            O => \N__13279\,
            I => \N__13276\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__13273\,
            I => ram_we_10
        );

    \I__1893\ : CEMux
    port map (
            O => \N__13270\,
            I => \N__13267\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__13267\,
            I => \N__13264\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__13264\,
            I => \N__13261\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__13261\,
            I => \N__13258\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__13258\,
            I => ram_we_8
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__13255\,
            I => \N__13251\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13243\
        );

    \I__1886\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13243\
        );

    \I__1885\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13243\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13240\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__13240\,
            I => \sb_translator_1.N_1088\
        );

    \I__1882\ : CEMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__1879\ : Sp12to4
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__13225\,
            I => ram_we_12
        );

    \I__1877\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13218\
        );

    \I__1876\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13215\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__13218\,
            I => \spi_slave_1.mosi_data_inZ0Z_5\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__13215\,
            I => \spi_slave_1.mosi_data_inZ0Z_5\
        );

    \I__1873\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13206\
        );

    \I__1872\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13203\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__13206\,
            I => \spi_slave_1.mosi_data_inZ0Z_6\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__13203\,
            I => \spi_slave_1.mosi_data_inZ0Z_6\
        );

    \I__1869\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13195\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13191\
        );

    \I__1867\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13188\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__13191\,
            I => \N__13185\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__13188\,
            I => \spi_slave_1.mosi_data_inZ0Z_7\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__13185\,
            I => \spi_slave_1.mosi_data_inZ0Z_7\
        );

    \I__1863\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13176\
        );

    \I__1862\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13173\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__13176\,
            I => \spi_slave_1.mosi_data_inZ0Z_4\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__13173\,
            I => \spi_slave_1.mosi_data_inZ0Z_4\
        );

    \I__1859\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13164\
        );

    \I__1858\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13161\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__13164\,
            I => \spi_slave_1.mosi_data_inZ0Z_0\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__13161\,
            I => \spi_slave_1.mosi_data_inZ0Z_0\
        );

    \I__1855\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13153\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__13153\,
            I => \N__13149\
        );

    \I__1853\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13146\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__13149\,
            I => \N__13138\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__13146\,
            I => \N__13138\
        );

    \I__1850\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13135\
        );

    \I__1849\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13132\
        );

    \I__1848\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13129\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__13138\,
            I => \N__13120\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13120\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__13132\,
            I => \N__13117\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__13129\,
            I => \N__13114\
        );

    \I__1843\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13111\
        );

    \I__1842\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13108\
        );

    \I__1841\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13104\
        );

    \I__1840\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13101\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__13120\,
            I => \N__13095\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__13117\,
            I => \N__13088\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__13114\,
            I => \N__13088\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13088\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__13108\,
            I => \N__13085\
        );

    \I__1834\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13082\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__13104\,
            I => \N__13077\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__13101\,
            I => \N__13077\
        );

    \I__1831\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13074\
        );

    \I__1830\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13071\
        );

    \I__1829\ : InMux
    port map (
            O => \N__13098\,
            I => \N__13067\
        );

    \I__1828\ : Span4Mux_s2_h
    port map (
            O => \N__13095\,
            I => \N__13062\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__13088\,
            I => \N__13062\
        );

    \I__1826\ : Span4Mux_s1_v
    port map (
            O => \N__13085\,
            I => \N__13057\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__13082\,
            I => \N__13057\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__13077\,
            I => \N__13050\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__13074\,
            I => \N__13050\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13050\
        );

    \I__1821\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13047\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__13067\,
            I => \N__13044\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__13062\,
            I => \N__13035\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__13057\,
            I => \N__13035\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__13050\,
            I => \N__13035\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13035\
        );

    \I__1815\ : Odrv12
    port map (
            O => \N__13044\,
            I => ram_data_in_0
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__13035\,
            I => ram_data_in_0
        );

    \I__1813\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13025\
        );

    \I__1812\ : InMux
    port map (
            O => \N__13029\,
            I => \N__13021\
        );

    \I__1811\ : InMux
    port map (
            O => \N__13028\,
            I => \N__13018\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__13025\,
            I => \N__13015\
        );

    \I__1809\ : InMux
    port map (
            O => \N__13024\,
            I => \N__13012\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__13021\,
            I => \N__13004\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__13018\,
            I => \N__13001\
        );

    \I__1806\ : Span4Mux_s1_v
    port map (
            O => \N__13015\,
            I => \N__12996\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__13012\,
            I => \N__12996\
        );

    \I__1804\ : InMux
    port map (
            O => \N__13011\,
            I => \N__12993\
        );

    \I__1803\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12990\
        );

    \I__1802\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12987\
        );

    \I__1801\ : InMux
    port map (
            O => \N__13008\,
            I => \N__12983\
        );

    \I__1800\ : InMux
    port map (
            O => \N__13007\,
            I => \N__12980\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__13004\,
            I => \N__12966\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__13001\,
            I => \N__12966\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__12996\,
            I => \N__12966\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__12993\,
            I => \N__12966\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__12990\,
            I => \N__12966\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12963\
        );

    \I__1793\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12960\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__12983\,
            I => \N__12955\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__12980\,
            I => \N__12955\
        );

    \I__1790\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12952\
        );

    \I__1789\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12949\
        );

    \I__1788\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12945\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__12966\,
            I => \N__12942\
        );

    \I__1786\ : Span4Mux_s1_v
    port map (
            O => \N__12963\,
            I => \N__12937\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12937\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__12955\,
            I => \N__12930\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__12952\,
            I => \N__12930\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__12949\,
            I => \N__12930\
        );

    \I__1781\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12927\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__12945\,
            I => \N__12924\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__12942\,
            I => \N__12915\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__12937\,
            I => \N__12915\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__12930\,
            I => \N__12915\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__12927\,
            I => \N__12915\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__12924\,
            I => ram_data_in_1
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__12915\,
            I => ram_data_in_1
        );

    \I__1773\ : InMux
    port map (
            O => \N__12910\,
            I => \N__12901\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12909\,
            I => \N__12898\
        );

    \I__1771\ : InMux
    port map (
            O => \N__12908\,
            I => \N__12891\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12888\
        );

    \I__1769\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12885\
        );

    \I__1768\ : InMux
    port map (
            O => \N__12905\,
            I => \N__12882\
        );

    \I__1767\ : InMux
    port map (
            O => \N__12904\,
            I => \N__12879\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__12901\,
            I => \N__12874\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__12898\,
            I => \N__12874\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12870\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12867\
        );

    \I__1762\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12863\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12894\,
            I => \N__12860\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__12891\,
            I => \N__12857\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__12888\,
            I => \N__12851\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__12885\,
            I => \N__12851\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__12882\,
            I => \N__12844\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12844\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__12874\,
            I => \N__12844\
        );

    \I__1754\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12841\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__12870\,
            I => \N__12838\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__12867\,
            I => \N__12835\
        );

    \I__1751\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12832\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__12863\,
            I => \N__12829\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12860\,
            I => \N__12824\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__12857\,
            I => \N__12824\
        );

    \I__1747\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12821\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__12851\,
            I => \N__12816\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__12844\,
            I => \N__12816\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__12841\,
            I => \N__12811\
        );

    \I__1743\ : Span4Mux_s1_v
    port map (
            O => \N__12838\,
            I => \N__12811\
        );

    \I__1742\ : Span4Mux_h
    port map (
            O => \N__12835\,
            I => \N__12808\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__12832\,
            I => \N__12801\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__12829\,
            I => \N__12801\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__12824\,
            I => \N__12801\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__12821\,
            I => \N__12796\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__12816\,
            I => \N__12796\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__12811\,
            I => \N__12789\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__12808\,
            I => \N__12789\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__12801\,
            I => \N__12789\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__12796\,
            I => ram_data_in_2
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__12789\,
            I => ram_data_in_2
        );

    \I__1731\ : InMux
    port map (
            O => \N__12784\,
            I => \N__12780\
        );

    \I__1730\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12772\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__12780\,
            I => \N__12768\
        );

    \I__1728\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12765\
        );

    \I__1727\ : InMux
    port map (
            O => \N__12778\,
            I => \N__12762\
        );

    \I__1726\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12758\
        );

    \I__1725\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12754\
        );

    \I__1724\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12748\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__12772\,
            I => \N__12745\
        );

    \I__1722\ : InMux
    port map (
            O => \N__12771\,
            I => \N__12742\
        );

    \I__1721\ : Span4Mux_h
    port map (
            O => \N__12768\,
            I => \N__12737\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__12765\,
            I => \N__12737\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__12762\,
            I => \N__12734\
        );

    \I__1718\ : InMux
    port map (
            O => \N__12761\,
            I => \N__12731\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__12758\,
            I => \N__12728\
        );

    \I__1716\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12725\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__12754\,
            I => \N__12722\
        );

    \I__1714\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12719\
        );

    \I__1713\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12716\
        );

    \I__1712\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12713\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__12748\,
            I => \N__12710\
        );

    \I__1710\ : Span4Mux_s1_v
    port map (
            O => \N__12745\,
            I => \N__12705\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__12742\,
            I => \N__12705\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__12737\,
            I => \N__12698\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__12734\,
            I => \N__12698\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__12731\,
            I => \N__12698\
        );

    \I__1705\ : Span4Mux_s1_v
    port map (
            O => \N__12728\,
            I => \N__12693\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__12725\,
            I => \N__12693\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__12722\,
            I => \N__12683\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__12719\,
            I => \N__12683\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__12716\,
            I => \N__12683\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12683\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__12710\,
            I => \N__12676\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__12705\,
            I => \N__12676\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__12698\,
            I => \N__12676\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__12693\,
            I => \N__12673\
        );

    \I__1695\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12670\
        );

    \I__1694\ : Span12Mux_s8_v
    port map (
            O => \N__12683\,
            I => \N__12665\
        );

    \I__1693\ : Sp12to4
    port map (
            O => \N__12676\,
            I => \N__12665\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__12673\,
            I => \N__12660\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12660\
        );

    \I__1690\ : Odrv12
    port map (
            O => \N__12665\,
            I => ram_data_in_3
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__12660\,
            I => ram_data_in_3
        );

    \I__1688\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12647\
        );

    \I__1687\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12644\
        );

    \I__1686\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12637\
        );

    \I__1685\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12632\
        );

    \I__1684\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12627\
        );

    \I__1683\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12624\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__12647\,
            I => \N__12619\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__12644\,
            I => \N__12619\
        );

    \I__1680\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12616\
        );

    \I__1679\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12613\
        );

    \I__1678\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12610\
        );

    \I__1677\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12607\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__12637\,
            I => \N__12604\
        );

    \I__1675\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12601\
        );

    \I__1674\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12598\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12595\
        );

    \I__1672\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12592\
        );

    \I__1671\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12589\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12584\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__12624\,
            I => \N__12584\
        );

    \I__1668\ : Span4Mux_s3_v
    port map (
            O => \N__12619\,
            I => \N__12577\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__12616\,
            I => \N__12577\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__12613\,
            I => \N__12577\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__12610\,
            I => \N__12574\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12569\
        );

    \I__1663\ : Span4Mux_s2_v
    port map (
            O => \N__12604\,
            I => \N__12569\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12566\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__12598\,
            I => \N__12561\
        );

    \I__1660\ : Span4Mux_s1_v
    port map (
            O => \N__12595\,
            I => \N__12561\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12554\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__12589\,
            I => \N__12554\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__12584\,
            I => \N__12554\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__12577\,
            I => \N__12547\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__12574\,
            I => \N__12547\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__12569\,
            I => \N__12547\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__12566\,
            I => \N__12540\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__12561\,
            I => \N__12540\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__12554\,
            I => \N__12540\
        );

    \I__1650\ : Span4Mux_h
    port map (
            O => \N__12547\,
            I => \N__12537\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__12540\,
            I => ram_data_in_4
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__12537\,
            I => ram_data_in_4
        );

    \I__1647\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12526\
        );

    \I__1646\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12526\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__1644\ : Span4Mux_h
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__12520\,
            I => mosi_data_out_8
        );

    \I__1642\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12514\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__12514\,
            I => \N__12509\
        );

    \I__1640\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12505\
        );

    \I__1639\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12502\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__12509\,
            I => \N__12499\
        );

    \I__1637\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12496\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__12505\,
            I => \N__12493\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__12502\,
            I => \sb_translator_1.cntZ0Z_0\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__12499\,
            I => \sb_translator_1.cntZ0Z_0\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__12496\,
            I => \sb_translator_1.cntZ0Z_0\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__12493\,
            I => \sb_translator_1.cntZ0Z_0\
        );

    \I__1631\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12478\
        );

    \I__1630\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12478\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__12475\,
            I => mosi_data_out_9
        );

    \I__1627\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12468\
        );

    \I__1626\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12465\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__12468\,
            I => \N__12462\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__12465\,
            I => \N__12458\
        );

    \I__1623\ : Span4Mux_h
    port map (
            O => \N__12462\,
            I => \N__12455\
        );

    \I__1622\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12452\
        );

    \I__1621\ : Span4Mux_s2_h
    port map (
            O => \N__12458\,
            I => \N__12449\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__12455\,
            I => \sb_translator_1.cntZ0Z_1\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__12452\,
            I => \sb_translator_1.cntZ0Z_1\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__12449\,
            I => \sb_translator_1.cntZ0Z_1\
        );

    \I__1617\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12439\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__12439\,
            I => \N__12435\
        );

    \I__1615\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12431\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__12435\,
            I => \N__12428\
        );

    \I__1613\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12425\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12422\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__12428\,
            I => \sb_translator_1.cntZ0Z_2\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__12425\,
            I => \sb_translator_1.cntZ0Z_2\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__12422\,
            I => \sb_translator_1.cntZ0Z_2\
        );

    \I__1608\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12409\
        );

    \I__1607\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12409\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__12409\,
            I => \N__12406\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__12406\,
            I => mosi_data_out_10
        );

    \I__1604\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12400\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__12400\,
            I => \N__12396\
        );

    \I__1602\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12393\
        );

    \I__1601\ : Odrv12
    port map (
            O => \N__12396\,
            I => \spi_slave_1.mosi_data_inZ0Z_16\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__12393\,
            I => \spi_slave_1.mosi_data_inZ0Z_16\
        );

    \I__1599\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12384\
        );

    \I__1598\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__12384\,
            I => \spi_slave_1.mosi_data_inZ0Z_3\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__12381\,
            I => \spi_slave_1.mosi_data_inZ0Z_3\
        );

    \I__1595\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12372\
        );

    \I__1594\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12369\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__12372\,
            I => \spi_slave_1.mosi_data_inZ0Z_2\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__12369\,
            I => \spi_slave_1.mosi_data_inZ0Z_2\
        );

    \I__1591\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12331\
        );

    \I__1590\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12331\
        );

    \I__1589\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12331\
        );

    \I__1588\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12331\
        );

    \I__1587\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12331\
        );

    \I__1586\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12331\
        );

    \I__1585\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12331\
        );

    \I__1584\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12331\
        );

    \I__1583\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12306\
        );

    \I__1582\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12306\
        );

    \I__1581\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12306\
        );

    \I__1580\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12306\
        );

    \I__1579\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12306\
        );

    \I__1578\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12306\
        );

    \I__1577\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12306\
        );

    \I__1576\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12306\
        );

    \I__1575\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12303\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__12331\,
            I => \N__12300\
        );

    \I__1573\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12283\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12283\
        );

    \I__1571\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12283\
        );

    \I__1570\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12283\
        );

    \I__1569\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12283\
        );

    \I__1568\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12283\
        );

    \I__1567\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12283\
        );

    \I__1566\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12283\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12278\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12278\
        );

    \I__1563\ : Span4Mux_h
    port map (
            O => \N__12300\,
            I => \N__12270\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__12283\,
            I => \N__12270\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__12278\,
            I => \N__12270\
        );

    \I__1560\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12264\
        );

    \I__1559\ : Sp12to4
    port map (
            O => \N__12270\,
            I => \N__12261\
        );

    \I__1558\ : InMux
    port map (
            O => \N__12269\,
            I => \N__12254\
        );

    \I__1557\ : InMux
    port map (
            O => \N__12268\,
            I => \N__12254\
        );

    \I__1556\ : InMux
    port map (
            O => \N__12267\,
            I => \N__12254\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__12264\,
            I => \spi_slave_1.clkZ0Z_0\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__12261\,
            I => \spi_slave_1.clkZ0Z_0\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__12254\,
            I => \spi_slave_1.clkZ0Z_0\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__12247\,
            I => \N__12241\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__12246\,
            I => \N__12237\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__12245\,
            I => \N__12233\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__12244\,
            I => \N__12229\
        );

    \I__1548\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12203\
        );

    \I__1547\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12203\
        );

    \I__1546\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12203\
        );

    \I__1545\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12203\
        );

    \I__1544\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12203\
        );

    \I__1543\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12203\
        );

    \I__1542\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12203\
        );

    \I__1541\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12203\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \N__12199\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12195\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12191\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__12224\,
            I => \N__12187\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \N__12183\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__12222\,
            I => \N__12179\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12175\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__12220\,
            I => \N__12171\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12167\
        );

    \I__1531\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12164\
        );

    \I__1530\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12147\
        );

    \I__1529\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12147\
        );

    \I__1528\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12147\
        );

    \I__1527\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12147\
        );

    \I__1526\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12147\
        );

    \I__1525\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12147\
        );

    \I__1524\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12147\
        );

    \I__1523\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12147\
        );

    \I__1522\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12129\
        );

    \I__1521\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12129\
        );

    \I__1520\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12129\
        );

    \I__1519\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12129\
        );

    \I__1518\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12129\
        );

    \I__1517\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12129\
        );

    \I__1516\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12129\
        );

    \I__1515\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12129\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__12167\,
            I => \N__12124\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__12164\,
            I => \N__12124\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12121\
        );

    \I__1511\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12118\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__12129\,
            I => \N__12113\
        );

    \I__1509\ : Sp12to4
    port map (
            O => \N__12124\,
            I => \N__12113\
        );

    \I__1508\ : Span12Mux_s3_v
    port map (
            O => \N__12121\,
            I => \N__12108\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__12118\,
            I => \N__12105\
        );

    \I__1506\ : Span12Mux_s10_v
    port map (
            O => \N__12113\,
            I => \N__12102\
        );

    \I__1505\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12097\
        );

    \I__1504\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12097\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__12108\,
            I => \spi_slave_1.clkZ0Z_1\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__12105\,
            I => \spi_slave_1.clkZ0Z_1\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__12102\,
            I => \spi_slave_1.clkZ0Z_1\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__12097\,
            I => \spi_slave_1.clkZ0Z_1\
        );

    \I__1499\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12084\
        );

    \I__1498\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12081\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__12084\,
            I => \N__12078\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__12081\,
            I => \N__12075\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__12078\,
            I => \N__12072\
        );

    \I__1494\ : Span4Mux_h
    port map (
            O => \N__12075\,
            I => \N__12069\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__12072\,
            I => \spi_slave_1.mosi_data_inZ0Z_17\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__12069\,
            I => \spi_slave_1.mosi_data_inZ0Z_17\
        );

    \I__1491\ : CEMux
    port map (
            O => \N__12064\,
            I => \N__12052\
        );

    \I__1490\ : CEMux
    port map (
            O => \N__12063\,
            I => \N__12052\
        );

    \I__1489\ : CEMux
    port map (
            O => \N__12062\,
            I => \N__12052\
        );

    \I__1488\ : CEMux
    port map (
            O => \N__12061\,
            I => \N__12052\
        );

    \I__1487\ : GlobalMux
    port map (
            O => \N__12052\,
            I => \N__12049\
        );

    \I__1486\ : gio2CtrlBuf
    port map (
            O => \N__12049\,
            I => \spi_slave_1.bitcnt_rxe_0_i_g\
        );

    \I__1485\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12042\
        );

    \I__1484\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12039\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__12042\,
            I => \N__12036\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12033\
        );

    \I__1481\ : Span4Mux_h
    port map (
            O => \N__12036\,
            I => \N__12030\
        );

    \I__1480\ : Span4Mux_h
    port map (
            O => \N__12033\,
            I => \N__12027\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__12030\,
            I => \spi_slave_1.mosi_data_inZ0Z_9\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__12027\,
            I => \spi_slave_1.mosi_data_inZ0Z_9\
        );

    \I__1477\ : InMux
    port map (
            O => \N__12022\,
            I => \N__12019\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__1475\ : Span4Mux_h
    port map (
            O => \N__12016\,
            I => \N__12012\
        );

    \I__1474\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12009\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__12012\,
            I => \spi_slave_1.mosi_data_inZ0Z_8\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__12009\,
            I => \spi_slave_1.mosi_data_inZ0Z_8\
        );

    \I__1471\ : InMux
    port map (
            O => \N__12004\,
            I => \N__12000\
        );

    \I__1470\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11997\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__12000\,
            I => \spi_slave_1.mosi_data_inZ0Z_10\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__11997\,
            I => \spi_slave_1.mosi_data_inZ0Z_10\
        );

    \I__1467\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11988\
        );

    \I__1466\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11985\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__11988\,
            I => \spi_slave_1.mosi_data_inZ0Z_11\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__11985\,
            I => \spi_slave_1.mosi_data_inZ0Z_11\
        );

    \I__1463\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11976\
        );

    \I__1462\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11973\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__11976\,
            I => \spi_slave_1.mosi_data_inZ0Z_12\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__11973\,
            I => \spi_slave_1.mosi_data_inZ0Z_12\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11964\
        );

    \I__1458\ : InMux
    port map (
            O => \N__11967\,
            I => \N__11961\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__11964\,
            I => \spi_slave_1.mosi_data_inZ0Z_13\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__11961\,
            I => \spi_slave_1.mosi_data_inZ0Z_13\
        );

    \I__1455\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11952\
        );

    \I__1454\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11949\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__11952\,
            I => \spi_slave_1.mosi_data_inZ0Z_14\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__11949\,
            I => \spi_slave_1.mosi_data_inZ0Z_14\
        );

    \I__1451\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11936\
        );

    \I__1450\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11936\
        );

    \I__1449\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11928\
        );

    \I__1448\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11928\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__11936\,
            I => \N__11925\
        );

    \I__1446\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11918\
        );

    \I__1445\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11918\
        );

    \I__1444\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11918\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__11928\,
            I => \spi_slave_1.bitcnt_txZ0Z_1\
        );

    \I__1442\ : Odrv12
    port map (
            O => \N__11925\,
            I => \spi_slave_1.bitcnt_txZ0Z_1\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__11918\,
            I => \spi_slave_1.bitcnt_txZ0Z_1\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__11911\,
            I => \spi_slave_1.m27_ns_1_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11905\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11902\
        );

    \I__1437\ : Span4Mux_s3_v
    port map (
            O => \N__11902\,
            I => \N__11899\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__11899\,
            I => \spi_slave_1.miso_RNOZ0Z_7\
        );

    \I__1435\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11893\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11890\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__11890\,
            I => \spi_slave_1.N_28_0\
        );

    \I__1432\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11884\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__11884\,
            I => \N__11881\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__11881\,
            I => \spi_slave_1.mosi_bufferZ0Z_1\
        );

    \I__1429\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11873\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__11877\,
            I => \N__11870\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__11876\,
            I => \N__11865\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11859\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11856\
        );

    \I__1424\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11851\
        );

    \I__1423\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11851\
        );

    \I__1422\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11848\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__11864\,
            I => \N__11845\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__11863\,
            I => \N__11842\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__11862\,
            I => \N__11838\
        );

    \I__1418\ : Span12Mux_s11_h
    port map (
            O => \N__11859\,
            I => \N__11835\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11832\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__11851\,
            I => \N__11829\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__11848\,
            I => \N__11826\
        );

    \I__1414\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11823\
        );

    \I__1413\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11820\
        );

    \I__1412\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11815\
        );

    \I__1411\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11815\
        );

    \I__1410\ : Span12Mux_v
    port map (
            O => \N__11835\,
            I => \N__11812\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__11832\,
            I => \N__11807\
        );

    \I__1408\ : Span4Mux_h
    port map (
            O => \N__11829\,
            I => \N__11807\
        );

    \I__1407\ : Span12Mux_s2_h
    port map (
            O => \N__11826\,
            I => \N__11798\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__11823\,
            I => \N__11798\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11798\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__11815\,
            I => \N__11798\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__11812\,
            I => cs_n
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__11807\,
            I => cs_n
        );

    \I__1401\ : Odrv12
    port map (
            O => \N__11798\,
            I => cs_n
        );

    \I__1400\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11788\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__1398\ : IoSpan4Mux
    port map (
            O => \N__11785\,
            I => \N__11782\
        );

    \I__1397\ : IoSpan4Mux
    port map (
            O => \N__11782\,
            I => \N__11779\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__11779\,
            I => mosi
        );

    \I__1395\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11773\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__11773\,
            I => \spi_slave_1.mosi_bufferZ0Z_0\
        );

    \I__1393\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11767\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__11767\,
            I => \N__11764\
        );

    \I__1391\ : Span4Mux_h
    port map (
            O => \N__11764\,
            I => \N__11761\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__11761\,
            I => \spi_slave_1.miso_data_outZ0Z_3\
        );

    \I__1389\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11755\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__11755\,
            I => \N__11752\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__11752\,
            I => \spi_slave_1.miso_data_outZ0Z_7\
        );

    \I__1386\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11746\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11743\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__11743\,
            I => \N__11740\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__11740\,
            I => miso_data_in_18
        );

    \I__1382\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11734\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__11734\,
            I => \spi_slave_1.miso_data_outZ0Z_2\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__11731\,
            I => \N__11728\
        );

    \I__1379\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11725\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__11725\,
            I => \spi_slave_1.miso_data_outZ0Z_18\
        );

    \I__1377\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__11719\,
            I => \N__11716\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__11716\,
            I => \N__11713\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__11713\,
            I => \spi_slave_1.m72_ns_1\
        );

    \I__1373\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11707\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__11707\,
            I => \spi_slave_1.miso_data_outZ0Z_14\
        );

    \I__1371\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__11701\,
            I => \spi_slave_1.miso_data_outZ0Z_13\
        );

    \I__1369\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11691\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__11697\,
            I => \N__11688\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__11696\,
            I => \N__11685\
        );

    \I__1366\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11680\
        );

    \I__1365\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11680\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__11691\,
            I => \N__11677\
        );

    \I__1363\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11672\
        );

    \I__1362\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11672\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__11680\,
            I => \spi_slave_1.bitcnt_txZ0Z_2\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__11677\,
            I => \spi_slave_1.bitcnt_txZ0Z_2\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__11672\,
            I => \spi_slave_1.bitcnt_txZ0Z_2\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \spi_slave_1.miso_RNOZ0Z_12_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__11653\,
            I => demux_data_in_55
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \demux.N_417_i_0_o2Z0Z_6_cascade_\
        );

    \I__1352\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11644\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__11644\,
            I => \demux.N_890\
        );

    \I__1350\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11638\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__11638\,
            I => demux_data_in_61
        );

    \I__1348\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11632\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__11629\,
            I => \N__11626\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__11626\,
            I => demux_data_in_77
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__11623\,
            I => \N__11620\
        );

    \I__1343\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__11617\,
            I => \N__11614\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__11614\,
            I => \N__11611\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__11611\,
            I => \N__11608\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__11608\,
            I => \N__11605\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__11605\,
            I => demux_data_in_85
        );

    \I__1337\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11599\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__1335\ : Span4Mux_h
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__1334\ : Span4Mux_s3_h
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__11590\,
            I => demux_data_in_53
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \demux.N_419_i_0_o2Z0Z_6_cascade_\
        );

    \I__1331\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11581\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__11581\,
            I => \demux.N_419_i_0_a3Z0Z_1\
        );

    \I__1329\ : InMux
    port map (
            O => \N__11578\,
            I => \N__11575\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__11575\,
            I => demux_data_in_60
        );

    \I__1327\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11569\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__11566\,
            I => \N__11563\
        );

    \I__1324\ : Span4Mux_h
    port map (
            O => \N__11563\,
            I => \N__11560\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__11560\,
            I => \N__11557\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__11557\,
            I => demux_data_in_84
        );

    \I__1321\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11551\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__11548\,
            I => \N__11545\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__11545\,
            I => demux_data_in_76
        );

    \I__1317\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11536\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__11536\,
            I => demux_data_in_52
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__11533\,
            I => \demux.N_420_i_0_o2Z0Z_6_cascade_\
        );

    \I__1313\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11527\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__11527\,
            I => \demux.N_420_i_0_a3Z0Z_1\
        );

    \I__1311\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11518\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__11518\,
            I => \N__11515\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__11515\,
            I => \spi_slave_1.miso_data_outZ0Z_6\
        );

    \I__1307\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__11506\,
            I => \spi_slave_1.miso_data_outZ0Z_1\
        );

    \I__1304\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__11500\,
            I => \N__11497\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__11497\,
            I => demux_data_in_54
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__11494\,
            I => \demux.N_877_cascade_\
        );

    \I__1300\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11488\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__11485\,
            I => demux_data_in_70
        );

    \I__1297\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__11479\,
            I => demux_data_in_62
        );

    \I__1295\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__11473\,
            I => \demux.N_418_i_0_o2Z0Z_6\
        );

    \I__1293\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__11455\,
            I => demux_data_in_83
        );

    \I__1287\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__11449\,
            I => demux_data_in_51
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__11446\,
            I => \demux.N_835_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11440\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__11440\,
            I => demux_data_in_59
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__1281\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11431\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__11428\,
            I => demux_data_in_67
        );

    \I__1278\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11422\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__11422\,
            I => \demux.N_421_i_0_o2Z0Z_6\
        );

    \I__1276\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__11416\,
            I => demux_data_in_63
        );

    \I__1274\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11410\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__11410\,
            I => demux_data_in_57
        );

    \I__1272\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11404\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11401\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__1269\ : Span4Mux_v
    port map (
            O => \N__11398\,
            I => \N__11395\
        );

    \I__1268\ : Span4Mux_h
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__11392\,
            I => demux_data_in_87
        );

    \I__1266\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11386\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__11386\,
            I => \N__11383\
        );

    \I__1264\ : Span4Mux_h
    port map (
            O => \N__11383\,
            I => \N__11380\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__11380\,
            I => demux_data_in_79
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__11377\,
            I => \N__11373\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__11376\,
            I => \N__11370\
        );

    \I__1260\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11362\
        );

    \I__1259\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11362\
        );

    \I__1258\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11362\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__11359\,
            I => \sb_translator_1.N_1092\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_\
        );

    \I__1254\ : CEMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__1252\ : Span4Mux_h
    port map (
            O => \N__11347\,
            I => \N__11344\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__11344\,
            I => \N__11341\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__11341\,
            I => ram_we_11
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__11338\,
            I => \sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_\
        );

    \I__1248\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11332\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__11332\,
            I => \N__11325\
        );

    \I__1246\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11316\
        );

    \I__1245\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11316\
        );

    \I__1244\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11316\
        );

    \I__1243\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11316\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__11325\,
            I => \N__11313\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11310\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__11313\,
            I => \N__11307\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__11310\,
            I => \N__11304\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__11307\,
            I => mosi_data_out_17
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__11304\,
            I => mosi_data_out_17
        );

    \I__1236\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11296\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__11284\,
            I => demux_data_in_86
        );

    \I__1230\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11275\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__11275\,
            I => \N__11271\
        );

    \I__1227\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11268\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__11271\,
            I => \N__11265\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11262\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__11265\,
            I => \N__11259\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__11262\,
            I => \N__11256\
        );

    \I__1222\ : Span4Mux_h
    port map (
            O => \N__11259\,
            I => \N__11253\
        );

    \I__1221\ : Span4Mux_h
    port map (
            O => \N__11256\,
            I => \N__11250\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__11253\,
            I => reset_n
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__11250\,
            I => reset_n
        );

    \I__1218\ : IoInMux
    port map (
            O => \N__11245\,
            I => \N__11242\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__11242\,
            I => \N__11239\
        );

    \I__1216\ : IoSpan4Mux
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__1215\ : Span4Mux_s3_v
    port map (
            O => \N__11236\,
            I => \N__11233\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__11233\,
            I => reset_n_i
        );

    \I__1213\ : CEMux
    port map (
            O => \N__11230\,
            I => \N__11227\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11224\
        );

    \I__1211\ : Span4Mux_s2_v
    port map (
            O => \N__11224\,
            I => \N__11221\
        );

    \I__1210\ : Span4Mux_h
    port map (
            O => \N__11221\,
            I => \N__11218\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__11218\,
            I => ram_we_3
        );

    \I__1208\ : CEMux
    port map (
            O => \N__11215\,
            I => \N__11212\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11209\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__11209\,
            I => \N__11206\
        );

    \I__1205\ : Span12Mux_s7_v
    port map (
            O => \N__11206\,
            I => \N__11203\
        );

    \I__1204\ : Odrv12
    port map (
            O => \N__11203\,
            I => ram_we_13
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_\
        );

    \I__1202\ : CEMux
    port map (
            O => \N__11197\,
            I => \N__11194\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__11194\,
            I => ram_we_5
        );

    \I__1200\ : CEMux
    port map (
            O => \N__11191\,
            I => \N__11188\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__11185\,
            I => \N__11182\
        );

    \I__1197\ : Span4Mux_s0_h
    port map (
            O => \N__11182\,
            I => \N__11179\
        );

    \I__1196\ : Span4Mux_h
    port map (
            O => \N__11179\,
            I => \N__11176\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__11176\,
            I => ram_we_7
        );

    \I__1194\ : CEMux
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11167\
        );

    \I__1192\ : Span12Mux_s7_v
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__11164\,
            I => ram_we_9
        );

    \I__1190\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11158\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11155\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__11155\,
            I => \N__11151\
        );

    \I__1187\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11148\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__11151\,
            I => \spi_slave_1.mosi_data_inZ0Z_1\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__11148\,
            I => \spi_slave_1.mosi_data_inZ0Z_1\
        );

    \I__1184\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11140\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__11140\,
            I => \N__11137\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__11137\,
            I => \sb_translator_1.un1_num_leds_n_9\
        );

    \I__1181\ : InMux
    port map (
            O => \N__11134\,
            I => \bfn_4_4_0_\
        );

    \I__1180\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11128\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11125\
        );

    \I__1178\ : Odrv12
    port map (
            O => \N__11125\,
            I => \sb_translator_1.un1_num_leds_n_10\
        );

    \I__1177\ : InMux
    port map (
            O => \N__11122\,
            I => \sb_translator_1.un1_num_leds_0_cry_9\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__11119\,
            I => \N__11116\
        );

    \I__1175\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11113\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11110\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__11110\,
            I => \sb_translator_1.un1_num_leds_n_11\
        );

    \I__1172\ : InMux
    port map (
            O => \N__11107\,
            I => \sb_translator_1.un1_num_leds_0_cry_10\
        );

    \I__1171\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11101\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__11101\,
            I => \N__11098\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__11098\,
            I => \sb_translator_1.un1_num_leds_n_12\
        );

    \I__1168\ : InMux
    port map (
            O => \N__11095\,
            I => \sb_translator_1.un1_num_leds_0_cry_11\
        );

    \I__1167\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11089\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__11089\,
            I => \N__11086\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__11086\,
            I => \sb_translator_1.un1_num_leds_n_13\
        );

    \I__1164\ : InMux
    port map (
            O => \N__11083\,
            I => \sb_translator_1.un1_num_leds_0_cry_12\
        );

    \I__1163\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11077\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__11077\,
            I => \N__11074\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__11074\,
            I => \sb_translator_1.un1_num_leds_n_14\
        );

    \I__1160\ : InMux
    port map (
            O => \N__11071\,
            I => \sb_translator_1.un1_num_leds_0_cry_13\
        );

    \I__1159\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11065\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__11065\,
            I => \N__11062\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__11062\,
            I => \sb_translator_1.un1_num_leds_n_15\
        );

    \I__1156\ : InMux
    port map (
            O => \N__11059\,
            I => \sb_translator_1.un1_num_leds_0_cry_14\
        );

    \I__1155\ : InMux
    port map (
            O => \N__11056\,
            I => \sb_translator_1.un1_num_leds_0_cry_15\
        );

    \I__1154\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11050\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__11050\,
            I => \N__11047\
        );

    \I__1152\ : Span4Mux_h
    port map (
            O => \N__11047\,
            I => \N__11044\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__11044\,
            I => \sb_translator_1.un1_num_leds_n_16\
        );

    \I__1150\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11038\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__11038\,
            I => \N__11035\
        );

    \I__1148\ : Odrv12
    port map (
            O => \N__11035\,
            I => \sb_translator_1.un1_num_leds_n_1\
        );

    \I__1147\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11029\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__11029\,
            I => \N__11026\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__11026\,
            I => \sb_translator_1.un1_num_leds_n_2\
        );

    \I__1144\ : InMux
    port map (
            O => \N__11023\,
            I => \sb_translator_1.un1_num_leds_0_cry_1\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__11020\,
            I => \N__11017\
        );

    \I__1142\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11014\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__11014\,
            I => \N__11011\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__11011\,
            I => \sb_translator_1.un1_num_leds_n_3\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11008\,
            I => \sb_translator_1.un1_num_leds_0_cry_2\
        );

    \I__1138\ : InMux
    port map (
            O => \N__11005\,
            I => \N__11002\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__11002\,
            I => \N__10999\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__10999\,
            I => \sb_translator_1.un1_num_leds_n_4\
        );

    \I__1135\ : InMux
    port map (
            O => \N__10996\,
            I => \sb_translator_1.un1_num_leds_0_cry_3\
        );

    \I__1134\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10990\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10987\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__10987\,
            I => \sb_translator_1.un1_num_leds_n_5\
        );

    \I__1131\ : InMux
    port map (
            O => \N__10984\,
            I => \sb_translator_1.un1_num_leds_0_cry_4\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__1129\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10975\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__10975\,
            I => \N__10972\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__10972\,
            I => \sb_translator_1.un1_num_leds_n_6\
        );

    \I__1126\ : InMux
    port map (
            O => \N__10969\,
            I => \sb_translator_1.un1_num_leds_0_cry_5\
        );

    \I__1125\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10963\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10960\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__10960\,
            I => \sb_translator_1.un1_num_leds_n_7\
        );

    \I__1122\ : InMux
    port map (
            O => \N__10957\,
            I => \sb_translator_1.un1_num_leds_0_cry_6\
        );

    \I__1121\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10951\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10948\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__10948\,
            I => \N__10945\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__10945\,
            I => \sb_translator_1.un1_num_leds_n_8\
        );

    \I__1117\ : InMux
    port map (
            O => \N__10942\,
            I => \sb_translator_1.un1_num_leds_0_cry_7\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__10939\,
            I => \spi_slave_1.N_49_0_cascade_\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__10936\,
            I => \spi_slave_1.N_25_0_cascade_\
        );

    \I__1114\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__10930\,
            I => \N__10927\
        );

    \I__1112\ : Span4Mux_s3_h
    port map (
            O => \N__10927\,
            I => \N__10924\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__10924\,
            I => \spi_slave_1.miso_data_outZ0Z_23\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__10921\,
            I => \N__10916\
        );

    \I__1109\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10911\
        );

    \I__1108\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10908\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10901\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10901\
        );

    \I__1105\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10901\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__10911\,
            I => \N__10898\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__10908\,
            I => \spi_slave_1.miso_data_out_0_sqmuxa\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__10901\,
            I => \spi_slave_1.miso_data_out_0_sqmuxa\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__10898\,
            I => \spi_slave_1.miso_data_out_0_sqmuxa\
        );

    \I__1100\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10888\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__10888\,
            I => \spi_slave_1.N_96_mux\
        );

    \I__1098\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10880\
        );

    \I__1097\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10877\
        );

    \I__1096\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10874\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__10880\,
            I => \spi_slave_1.N_94_mux\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__10877\,
            I => \spi_slave_1.N_94_mux\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__10874\,
            I => \spi_slave_1.N_94_mux\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10867\,
            I => \spi_slave_1.N_94_mux_cascade_\
        );

    \I__1091\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10852\
        );

    \I__1090\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10852\
        );

    \I__1089\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10852\
        );

    \I__1088\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10849\
        );

    \I__1087\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10846\
        );

    \I__1086\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10843\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10852\,
            I => \N__10840\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__10849\,
            I => \spi_slave_1.bitcnt_txZ0Z_3\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__10846\,
            I => \spi_slave_1.bitcnt_txZ0Z_3\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__10843\,
            I => \spi_slave_1.bitcnt_txZ0Z_3\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__10840\,
            I => \spi_slave_1.bitcnt_txZ0Z_3\
        );

    \I__1080\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10825\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10825\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__10825\,
            I => \spi_slave_1.N_17_0\
        );

    \I__1077\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10819\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__10819\,
            I => \spi_slave_1.N_20_0\
        );

    \I__1075\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10813\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__10813\,
            I => \spi_slave_1.N_91\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__10810\,
            I => \N__10807\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10807\,
            I => \N__10803\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10800\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__10803\,
            I => miso
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__10800\,
            I => miso
        );

    \I__1068\ : IoInMux
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10789\
        );

    \I__1066\ : IoSpan4Mux
    port map (
            O => \N__10789\,
            I => \N__10786\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__10786\,
            I => \spi_slave_1.bitcnt_rxe_0_i\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__10783\,
            I => \N__10780\
        );

    \I__1063\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__10777\,
            I => \spi_slave_1.bitcnt_tx10\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__10774\,
            I => \spi_slave_1.bitcnt_tx10_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10768\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__10768\,
            I => \N__10765\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__10765\,
            I => \spi_slave_1.miso_data_outZ0Z_8\
        );

    \I__1057\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10758\
        );

    \I__1056\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__10755\,
            I => \N__10747\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__10752\,
            I => \N__10747\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__10747\,
            I => miso_tx
        );

    \I__1051\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10741\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__10741\,
            I => \N__10738\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__10738\,
            I => \spi_slave_1.N_82\
        );

    \I__1048\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10732\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__10732\,
            I => \spi_slave_1.miso_RNOZ0Z_17\
        );

    \I__1046\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10726\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__10723\,
            I => \spi_slave_1.miso_RNOZ0Z_10\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__10720\,
            I => \spi_slave_1.m48_ns_1_cascade_\
        );

    \I__1042\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10714\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__10714\,
            I => miso_data_in_8
        );

    \I__1040\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__1039\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10705\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__10705\,
            I => \N__10699\
        );

    \I__1037\ : InMux
    port map (
            O => \N__10704\,
            I => \N__10692\
        );

    \I__1036\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10692\
        );

    \I__1035\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10692\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__10699\,
            I => \spi_slave_1.clk_pos_i\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__10692\,
            I => \spi_slave_1.clk_pos_i\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__10687\,
            I => \N__10684\
        );

    \I__1031\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10681\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__10681\,
            I => \spi_slave_1.miso_data_outZ0Z_22\
        );

    \I__1029\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10675\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__10675\,
            I => \spi_slave_1.miso_data_outZ0Z_21\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__10672\,
            I => \spi_slave_1.m81_ns_1_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10666\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__10666\,
            I => \spi_slave_1.miso_data_outZ0Z_5\
        );

    \I__1024\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10660\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__10660\,
            I => \spi_slave_1.miso_data_outZ0Z_4\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__10657\,
            I => \N__10654\
        );

    \I__1021\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10651\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__10651\,
            I => \spi_slave_1.miso_data_outZ0Z_20\
        );

    \I__1019\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10645\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__10645\,
            I => \spi_slave_1.miso_data_outZ0Z_19\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__10642\,
            I => \spi_slave_1.m60_ns_1_cascade_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10636\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__10636\,
            I => \N__10633\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__10633\,
            I => clk_spi
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__10630\,
            I => \N__10626\
        );

    \I__1012\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10623\
        );

    \I__1011\ : InMux
    port map (
            O => \N__10626\,
            I => \N__10620\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__10623\,
            I => \sb_translator_1.instr_tmpZ0Z_22\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__10620\,
            I => \sb_translator_1.instr_tmpZ0Z_22\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__10615\,
            I => \N__10611\
        );

    \I__1007\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10608\
        );

    \I__1006\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10605\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__10608\,
            I => \sb_translator_1.instr_tmpZ0Z_23\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__10605\,
            I => \sb_translator_1.instr_tmpZ0Z_23\
        );

    \I__1003\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10597\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__10597\,
            I => miso_data_in_19
        );

    \I__1001\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10591\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__10591\,
            I => miso_data_in_20
        );

    \I__999\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10585\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__10585\,
            I => miso_data_in_21
        );

    \I__997\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10579\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__10579\,
            I => miso_data_in_22
        );

    \I__995\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10573\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__10573\,
            I => miso_data_in_23
        );

    \I__993\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10567\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__10567\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_9\
        );

    \I__991\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10561\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10553\
        );

    \I__989\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10544\
        );

    \I__988\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10544\
        );

    \I__987\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10544\
        );

    \I__986\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10544\
        );

    \I__985\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10541\
        );

    \I__984\ : Span4Mux_s2_h
    port map (
            O => \N__10553\,
            I => \N__10538\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__10544\,
            I => \sb_translator_1.cntZ0Z_9\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__10541\,
            I => \sb_translator_1.cntZ0Z_9\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__10538\,
            I => \sb_translator_1.cntZ0Z_9\
        );

    \I__980\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10526\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__10530\,
            I => \N__10523\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__10529\,
            I => \N__10519\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__10526\,
            I => \N__10514\
        );

    \I__976\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10505\
        );

    \I__975\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10505\
        );

    \I__974\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10505\
        );

    \I__973\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10505\
        );

    \I__972\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10502\
        );

    \I__971\ : Span4Mux_s2_h
    port map (
            O => \N__10514\,
            I => \N__10499\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__10505\,
            I => \sb_translator_1.cntZ0Z_12\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__10502\,
            I => \sb_translator_1.cntZ0Z_12\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__10499\,
            I => \sb_translator_1.cntZ0Z_12\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__10492\,
            I => \N__10488\
        );

    \I__966\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10485\
        );

    \I__965\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10482\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__10485\,
            I => \sb_translator_1.instr_tmpZ0Z_18\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__10482\,
            I => \sb_translator_1.instr_tmpZ0Z_18\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__10477\,
            I => \N__10473\
        );

    \I__961\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10470\
        );

    \I__960\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10467\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__10470\,
            I => \sb_translator_1.instr_tmpZ0Z_19\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__10467\,
            I => \sb_translator_1.instr_tmpZ0Z_19\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__10462\,
            I => \N__10458\
        );

    \I__956\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10455\
        );

    \I__955\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10452\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__10455\,
            I => \sb_translator_1.instr_tmpZ0Z_20\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__10452\,
            I => \sb_translator_1.instr_tmpZ0Z_20\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__10447\,
            I => \N__10443\
        );

    \I__951\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10440\
        );

    \I__950\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10437\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__10440\,
            I => \sb_translator_1.instr_tmpZ0Z_21\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__10437\,
            I => \sb_translator_1.instr_tmpZ0Z_21\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__10432\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_0_cascade_\
        );

    \I__946\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10426\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__10426\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_13\
        );

    \I__944\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10419\
        );

    \I__943\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10416\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__10419\,
            I => \N__10413\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__10416\,
            I => \sb_translator_1.cntZ0Z_13\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__10413\,
            I => \sb_translator_1.cntZ0Z_13\
        );

    \I__939\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10405\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__10405\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_14\
        );

    \I__937\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10398\
        );

    \I__936\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10395\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__10398\,
            I => \N__10392\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__10395\,
            I => \sb_translator_1.cntZ0Z_14\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__10392\,
            I => \sb_translator_1.cntZ0Z_14\
        );

    \I__932\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10384\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__10384\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_15\
        );

    \I__930\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10377\
        );

    \I__929\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10374\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__10377\,
            I => \N__10371\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__10374\,
            I => \sb_translator_1.cntZ0Z_15\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__10371\,
            I => \sb_translator_1.cntZ0Z_15\
        );

    \I__925\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10363\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__10363\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_16\
        );

    \I__923\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10356\
        );

    \I__922\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10353\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__10356\,
            I => \sb_translator_1.cntZ0Z_16\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__10353\,
            I => \sb_translator_1.cntZ0Z_16\
        );

    \I__919\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10345\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__10345\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_1\
        );

    \I__917\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10339\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__10339\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_11\
        );

    \I__915\ : InMux
    port map (
            O => \N__10336\,
            I => \N__10333\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__10333\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_12\
        );

    \I__913\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10327\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__10327\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_10\
        );

    \I__911\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10321\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__10321\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_2\
        );

    \I__909\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__10315\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_3\
        );

    \I__907\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10309\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__10309\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_4\
        );

    \I__905\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10303\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__10303\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_5\
        );

    \I__903\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10297\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__10297\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_6\
        );

    \I__901\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__10291\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_7\
        );

    \I__899\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__10285\,
            I => \sb_translator_1.cnt_RNO_0Z0Z_8\
        );

    \I__897\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10278\
        );

    \I__896\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10275\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__10278\,
            I => \sb_translator_1.stateZ0Z_5\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__10275\,
            I => \sb_translator_1.stateZ0Z_5\
        );

    \I__893\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10267\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__10267\,
            I => \spi_slave_1.mosi_data_inZ0Z_23\
        );

    \I__891\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10260\
        );

    \I__890\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__10260\,
            I => \spi_slave_1.mosi_data_inZ0Z_18\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__10257\,
            I => \spi_slave_1.mosi_data_inZ0Z_18\
        );

    \I__887\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10248\
        );

    \I__886\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10245\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__10248\,
            I => \spi_slave_1.mosi_data_inZ0Z_19\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__10245\,
            I => \spi_slave_1.mosi_data_inZ0Z_19\
        );

    \I__883\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10236\
        );

    \I__882\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10233\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__10236\,
            I => \spi_slave_1.mosi_data_inZ0Z_20\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__10233\,
            I => \spi_slave_1.mosi_data_inZ0Z_20\
        );

    \I__879\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10224\
        );

    \I__878\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10221\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__10224\,
            I => \spi_slave_1.mosi_data_inZ0Z_21\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__10221\,
            I => \spi_slave_1.mosi_data_inZ0Z_21\
        );

    \I__875\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10212\
        );

    \I__874\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10209\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__10212\,
            I => \spi_slave_1.mosi_data_inZ0Z_22\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__10209\,
            I => \spi_slave_1.mosi_data_inZ0Z_22\
        );

    \I__871\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10201\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__10201\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO\
        );

    \I__869\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__10195\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO\
        );

    \I__867\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10188\
        );

    \I__866\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10185\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__10188\,
            I => \spi_slave_1.bitcnt_rxZ0Z_3\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__10185\,
            I => \spi_slave_1.bitcnt_rxZ0Z_3\
        );

    \I__863\ : InMux
    port map (
            O => \N__10180\,
            I => \spi_slave_1.bitcnt_rx_cry_2\
        );

    \I__862\ : InMux
    port map (
            O => \N__10177\,
            I => \spi_slave_1.bitcnt_rx_cry_3\
        );

    \I__861\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10169\
        );

    \I__860\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10164\
        );

    \I__859\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10164\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__10169\,
            I => \spi_slave_1.bitcnt_rxZ0Z_4\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__10164\,
            I => \spi_slave_1.bitcnt_rxZ0Z_4\
        );

    \I__856\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10156\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__10156\,
            I => miso_en
        );

    \I__854\ : InMux
    port map (
            O => \N__10153\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__10150\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_1\
        );

    \I__852\ : InMux
    port map (
            O => \N__10147\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_2\
        );

    \I__851\ : InMux
    port map (
            O => \N__10144\,
            I => \spi_slave_1.un1_bitcnt_tx_1_cry_3\
        );

    \I__850\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10138\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__10138\,
            I => \spi_slave_1.un3_mosi_data_out_3\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__10135\,
            I => \spi_slave_1.un3_mosi_data_out_3_cascade_\
        );

    \I__847\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10127\
        );

    \I__846\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10122\
        );

    \I__845\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10122\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__10127\,
            I => \spi_slave_1.bitcnt_rxZ0Z_0\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__10122\,
            I => \spi_slave_1.bitcnt_rxZ0Z_0\
        );

    \I__842\ : InMux
    port map (
            O => \N__10117\,
            I => \bfn_1_10_0_\
        );

    \I__841\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10110\
        );

    \I__840\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__10110\,
            I => \spi_slave_1.bitcnt_rxZ0Z_1\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__10107\,
            I => \spi_slave_1.bitcnt_rxZ0Z_1\
        );

    \I__837\ : InMux
    port map (
            O => \N__10102\,
            I => \spi_slave_1.bitcnt_rx_cry_0\
        );

    \I__836\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10095\
        );

    \I__835\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10092\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__10095\,
            I => \spi_slave_1.bitcnt_rxZ0Z_2\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__10092\,
            I => \spi_slave_1.bitcnt_rxZ0Z_2\
        );

    \I__832\ : InMux
    port map (
            O => \N__10087\,
            I => \spi_slave_1.bitcnt_rx_cry_1\
        );

    \I__831\ : InMux
    port map (
            O => \N__10084\,
            I => \sb_translator_1.cnt19_cry_31\
        );

    \I__830\ : InMux
    port map (
            O => \N__10081\,
            I => \sb_translator_1.cnt19_cry_32\
        );

    \I__829\ : InMux
    port map (
            O => \N__10078\,
            I => \bfn_1_7_0_\
        );

    \I__828\ : InMux
    port map (
            O => \N__10075\,
            I => \sb_translator_1.cnt19_cry_34\
        );

    \I__827\ : InMux
    port map (
            O => \N__10072\,
            I => \sb_translator_1.cnt19_cry_35\
        );

    \I__826\ : IoInMux
    port map (
            O => \N__10069\,
            I => \N__10066\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10063\
        );

    \I__824\ : Span4Mux_s1_v
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__10057\,
            I => \spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4\
        );

    \I__821\ : InMux
    port map (
            O => \N__10054\,
            I => \sb_translator_1.cnt19_cry_22\
        );

    \I__820\ : InMux
    port map (
            O => \N__10051\,
            I => \sb_translator_1.cnt19_cry_23\
        );

    \I__819\ : InMux
    port map (
            O => \N__10048\,
            I => \sb_translator_1.cnt19_cry_24\
        );

    \I__818\ : InMux
    port map (
            O => \N__10045\,
            I => \bfn_1_6_0_\
        );

    \I__817\ : InMux
    port map (
            O => \N__10042\,
            I => \sb_translator_1.cnt19_cry_26\
        );

    \I__816\ : InMux
    port map (
            O => \N__10039\,
            I => \sb_translator_1.cnt19_cry_27\
        );

    \I__815\ : InMux
    port map (
            O => \N__10036\,
            I => \sb_translator_1.cnt19_cry_28\
        );

    \I__814\ : InMux
    port map (
            O => \N__10033\,
            I => \sb_translator_1.cnt19_cry_29\
        );

    \I__813\ : InMux
    port map (
            O => \N__10030\,
            I => \sb_translator_1.cnt19_cry_30\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__10027\,
            I => \N__10024\
        );

    \I__811\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10021\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__10021\,
            I => \N__10018\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__10018\,
            I => \sb_translator_1.cnt_RNI0G0QZ0Z_13\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__10015\,
            I => \N__10012\
        );

    \I__807\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10009\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__10006\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__10006\,
            I => \sb_translator_1.cnt_RNI4L1QZ0Z_14\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__10003\,
            I => \N__10000\
        );

    \I__803\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9997\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__9997\,
            I => \N__9994\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__9994\,
            I => \sb_translator_1.cnt_RNI8Q2QZ0Z_15\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__9991\,
            I => \N__9988\
        );

    \I__799\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9985\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__9985\,
            I => \sb_translator_1.cnt_i_16\
        );

    \I__797\ : InMux
    port map (
            O => \N__9982\,
            I => \sb_translator_1.cnt19_cry_16\
        );

    \I__796\ : InMux
    port map (
            O => \N__9979\,
            I => \sb_translator_1.cnt19_cry_18\
        );

    \I__795\ : InMux
    port map (
            O => \N__9976\,
            I => \sb_translator_1.cnt19_cry_20\
        );

    \I__794\ : InMux
    port map (
            O => \N__9973\,
            I => \sb_translator_1.cnt19_cry_21\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__9970\,
            I => \N__9967\
        );

    \I__792\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9964\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__9964\,
            I => \sb_translator_1.cnt_RNI0T5OZ0Z_4\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__9961\,
            I => \N__9958\
        );

    \I__789\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9955\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__9955\,
            I => \sb_translator_1.cnt_RNI427OZ0Z_5\
        );

    \I__787\ : InMux
    port map (
            O => \N__9952\,
            I => \N__9949\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__9949\,
            I => \sb_translator_1.cnt_RNI878OZ0Z_6\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__9946\,
            I => \N__9943\
        );

    \I__784\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9940\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__9940\,
            I => \sb_translator_1.cnt_RNICC9OZ0Z_7\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \N__9934\
        );

    \I__781\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__9931\,
            I => \sb_translator_1.cnt_RNIGHAOZ0Z_8\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__9928\,
            I => \N__9925\
        );

    \I__778\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__9922\,
            I => \sb_translator_1.cnt_RNIKMBOZ0Z_9\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__9919\,
            I => \N__9916\
        );

    \I__775\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9913\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__9913\,
            I => \sb_translator_1.cnt_RNI6O3VZ0Z_10\
        );

    \I__773\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__9907\,
            I => \sb_translator_1.cnt_RNIO5UPZ0Z_11\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__9904\,
            I => \N__9901\
        );

    \I__770\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__9898\,
            I => \sb_translator_1.cnt_RNISAVPZ0Z_12\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__9895\,
            I => \N__9892\
        );

    \I__767\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9889\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__9889\,
            I => \sb_translator_1.cnt_i_0\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__9886\,
            I => \N__9883\
        );

    \I__764\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9880\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__9880\,
            I => \sb_translator_1.cnt_i_1\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__9877\,
            I => \N__9874\
        );

    \I__761\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9871\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__9871\,
            I => \sb_translator_1.cnt_RNIOI3OZ0Z_2\
        );

    \I__759\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9865\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__9865\,
            I => \sb_translator_1.cnt_RNISN4OZ0Z_3\
        );

    \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27512\
        );

    \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27519\
        );

    \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27462\
        );

    \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27430\
        );

    \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27477\
        );

    \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27446\
        );

    \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27423\
        );

    \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27442\
        );

    \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27419\
        );

    \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27504\
        );

    \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27491\
        );

    \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27456\
        );

    \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27472\
        );

    \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN\ : INV
    port map (
            O => \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net\,
            I => \N__27487\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.state56_a_5_cry_6\,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.state56_a_5_cry_14\,
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ws2812.un6_data_cry_7\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ws2812.un1_bit_counter_12_cry_7\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.un1_num_leds_0_cry_8\,
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt_leds_cry_7\,
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt_leds_cry_15\,
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt19_cry_7\,
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt19_cry_15\,
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt19_cry_25\,
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sb_translator_1.cnt19_cry_33\,
            carryinitout => \bfn_1_7_0_\
        );

    \sb_translator_1.state_RNI6JH4_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22798\,
            GLOBALBUFFEROUTPUT => \sb_translator_1.state_g_1\
        );

    \OSCInst0\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b00"
        )
    port map (
            CLKHFPU => \N__26124\,
            CLKHFEN => \N__26123\,
            CLKHF => clk_sb
        );

    \sb_translator_1.state_leds_RNIVONR_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18010\,
            GLOBALBUFFEROUTPUT => \sb_translator_1.state_leds_2_sqmuxa_g\
        );

    \reset_n_input_RNIVGR4_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11245\,
            GLOBALBUFFEROUTPUT => reset_n_i_g
        );

    \spi_slave_1.bitcnt_rx_RNIPNM61_0_4\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10069\,
            GLOBALBUFFEROUTPUT => \spi_slave_1.un3_mosi_data_out_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \spi_slave_1.clk_RNIVAC01_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10795\,
            GLOBALBUFFEROUTPUT => \spi_slave_1.bitcnt_rxe_0_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \sb_translator_1.instr_tx_LC_0_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__23998\,
            in1 => \N__10761\,
            in2 => \_gnd_net_\,
            in3 => \N__22072\,
            lcout => miso_tx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27439\,
            ce => 'H',
            sr => \N__27107\
        );

    \sb_translator_1.cnt_RNI4OM7_0_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12513\,
            in1 => \N__19108\,
            in2 => \N__9895\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_i_0\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \sb_translator_1.cnt19_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI1TPB_1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11041\,
            in2 => \N__9886\,
            in3 => \N__12471\,
            lcout => \sb_translator_1.cnt_i_1\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_0\,
            carryout => \sb_translator_1.cnt19_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIOI3O_2_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11032\,
            in2 => \N__9877\,
            in3 => \N__12438\,
            lcout => \sb_translator_1.cnt_RNIOI3OZ0Z_2\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_1\,
            carryout => \sb_translator_1.cnt19_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNISN4O_3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9868\,
            in2 => \N__11020\,
            in3 => \N__14628\,
            lcout => \sb_translator_1.cnt_RNISN4OZ0Z_3\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_2\,
            carryout => \sb_translator_1.cnt19_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI0T5O_4_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11005\,
            in2 => \N__9970\,
            in3 => \N__22560\,
            lcout => \sb_translator_1.cnt_RNI0T5OZ0Z_4\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_3\,
            carryout => \sb_translator_1.cnt19_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI427O_5_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10993\,
            in2 => \N__9961\,
            in3 => \N__14589\,
            lcout => \sb_translator_1.cnt_RNI427OZ0Z_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_4\,
            carryout => \sb_translator_1.cnt19_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI878O_6_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22506\,
            in1 => \N__9952\,
            in2 => \N__10981\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_RNI878OZ0Z_6\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_5\,
            carryout => \sb_translator_1.cnt19_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNICC9O_7_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10966\,
            in2 => \N__9946\,
            in3 => \N__22927\,
            lcout => \sb_translator_1.cnt_RNICC9OZ0Z_7\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_6\,
            carryout => \sb_translator_1.cnt19_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIGHAO_8_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10954\,
            in2 => \N__9937\,
            in3 => \N__21446\,
            lcout => \sb_translator_1.cnt_RNIGHAOZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => \sb_translator_1.cnt19_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIKMBO_9_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11143\,
            in2 => \N__9928\,
            in3 => \N__10564\,
            lcout => \sb_translator_1.cnt_RNIKMBOZ0Z_9\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_8\,
            carryout => \sb_translator_1.cnt19_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI6O3V_10_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11131\,
            in2 => \N__9919\,
            in3 => \N__17291\,
            lcout => \sb_translator_1.cnt_RNI6O3VZ0Z_10\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_9\,
            carryout => \sb_translator_1.cnt19_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIO5UP_11_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17358\,
            in1 => \N__9910\,
            in2 => \N__11119\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_RNIO5UPZ0Z_11\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_10\,
            carryout => \sb_translator_1.cnt19_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNISAVP_12_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11104\,
            in2 => \N__9904\,
            in3 => \N__10531\,
            lcout => \sb_translator_1.cnt_RNISAVPZ0Z_12\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_11\,
            carryout => \sb_translator_1.cnt19_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI0G0Q_13_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11092\,
            in2 => \N__10027\,
            in3 => \N__10423\,
            lcout => \sb_translator_1.cnt_RNI0G0QZ0Z_13\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_12\,
            carryout => \sb_translator_1.cnt19_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI4L1Q_14_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10402\,
            in1 => \N__11080\,
            in2 => \N__10015\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_RNI4L1QZ0Z_14\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_13\,
            carryout => \sb_translator_1.cnt19_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNI8Q2Q_15_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11068\,
            in2 => \N__10003\,
            in3 => \N__10381\,
            lcout => \sb_translator_1.cnt_RNI8Q2QZ0Z_15\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_14\,
            carryout => \sb_translator_1.cnt19_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIQ4UI_16_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11053\,
            in2 => \N__9991\,
            in3 => \N__10359\,
            lcout => \sb_translator_1.cnt_i_16\,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \sb_translator_1.cnt19_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNIOCIR9_5_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__10281\,
            in1 => \N__23011\,
            in2 => \_gnd_net_\,
            in3 => \N__9982\,
            lcout => \sb_translator_1.state_RNIOCIR9Z0Z_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_16\,
            carryout => \sb_translator_1.cnt19_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt19_cry_18_THRU_LUT4_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12508\,
            in2 => \_gnd_net_\,
            in3 => \N__9979\,
            lcout => \sb_translator_1.cnt19_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_18\,
            carryout => \sb_translator_1.cnt19_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_1_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12461\,
            in2 => \_gnd_net_\,
            in3 => \N__9976\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_20\,
            carryout => \sb_translator_1.cnt19_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_2_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12434\,
            in2 => \_gnd_net_\,
            in3 => \N__9973\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_21\,
            carryout => \sb_translator_1.cnt19_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_3_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14624\,
            in2 => \_gnd_net_\,
            in3 => \N__10054\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_22\,
            carryout => \sb_translator_1.cnt19_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_4_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22556\,
            in2 => \_gnd_net_\,
            in3 => \N__10051\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_23\,
            carryout => \sb_translator_1.cnt19_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_5_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14585\,
            in2 => \_gnd_net_\,
            in3 => \N__10048\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_24\,
            carryout => \sb_translator_1.cnt19_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_6_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22502\,
            in2 => \_gnd_net_\,
            in3 => \N__10045\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \sb_translator_1.cnt19_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_7_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22919\,
            in2 => \_gnd_net_\,
            in3 => \N__10042\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_26\,
            carryout => \sb_translator_1.cnt19_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_8_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21447\,
            in2 => \_gnd_net_\,
            in3 => \N__10039\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_27\,
            carryout => \sb_translator_1.cnt19_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_9_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10556\,
            in2 => \_gnd_net_\,
            in3 => \N__10036\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_28\,
            carryout => \sb_translator_1.cnt19_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_10_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17292\,
            in2 => \_gnd_net_\,
            in3 => \N__10033\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_29\,
            carryout => \sb_translator_1.cnt19_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_11_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17346\,
            in2 => \_gnd_net_\,
            in3 => \N__10030\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_30\,
            carryout => \sb_translator_1.cnt19_cry_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_12_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10517\,
            in2 => \_gnd_net_\,
            in3 => \N__10084\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_31\,
            carryout => \sb_translator_1.cnt19_cry_32\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_13_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10422\,
            in2 => \_gnd_net_\,
            in3 => \N__10081\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_32\,
            carryout => \sb_translator_1.cnt19_cry_33\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_14_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10401\,
            in2 => \_gnd_net_\,
            in3 => \N__10078\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \sb_translator_1.cnt19_cry_34\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_15_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10380\,
            in2 => \_gnd_net_\,
            in3 => \N__10075\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt19_cry_34\,
            carryout => \sb_translator_1.cnt19_cry_35\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNO_0_16_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10360\,
            in2 => \_gnd_net_\,
            in3 => \N__10072\,
            lcout => \sb_translator_1.cnt_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNIKJOC_5_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__10282\,
            in1 => \N__22066\,
            in2 => \_gnd_net_\,
            in3 => \N__16853\,
            lcout => \sb_translator_1.state_RNIKJOCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_tmp_23_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__16844\,
            in1 => \N__22762\,
            in2 => \N__10615\,
            in3 => \N__22071\,
            lcout => \sb_translator_1.instr_tmpZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27434\,
            ce => 'H',
            sr => \N__27088\
        );

    \sb_translator_1.instr_tmp_21_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__16843\,
            in1 => \N__22070\,
            in2 => \N__10447\,
            in3 => \N__22644\,
            lcout => \sb_translator_1.instr_tmpZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27434\,
            ce => 'H',
            sr => \N__27088\
        );

    \sb_translator_1.instr_tmp_18_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17680\,
            in1 => \N__22073\,
            in2 => \N__10492\,
            in3 => \N__16842\,
            lcout => \sb_translator_1.instr_tmpZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27434\,
            ce => 'H',
            sr => \N__27088\
        );

    \spi_slave_1.bitcnt_rx_RNIPNM61_4_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10172\,
            in1 => \N__10141\,
            in2 => \_gnd_net_\,
            in3 => \N__10130\,
            lcout => \spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_rx_RNI3EGR_1_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10191\,
            in1 => \N__10098\,
            in2 => \N__11876\,
            in3 => \N__10113\,
            lcout => \spi_slave_1.un3_mosi_data_out_3\,
            ltout => \spi_slave_1.un3_mosi_data_out_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.mosi_rx_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__10173\,
            in1 => \_gnd_net_\,
            in2 => \N__10135\,
            in3 => \N__10131\,
            lcout => mosi_rx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27440\,
            ce => 'H',
            sr => \N__27095\
        );

    \sb_translator_1.instr_tmp_19_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__22064\,
            in1 => \N__17623\,
            in2 => \N__10477\,
            in3 => \N__16826\,
            lcout => \sb_translator_1.instr_tmpZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27440\,
            ce => 'H',
            sr => \N__27095\
        );

    \sb_translator_1.instr_tmp_20_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__16827\,
            in1 => \N__17572\,
            in2 => \N__10462\,
            in3 => \N__22065\,
            lcout => \sb_translator_1.instr_tmpZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27440\,
            ce => 'H',
            sr => \N__27095\
        );

    \sb_translator_1.state_RNIH20C_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22063\,
            in1 => \N__16825\,
            in2 => \_gnd_net_\,
            in3 => \N__22643\,
            lcout => \sb_translator_1.N_1087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_6_0_0_a2_1_9_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17622\,
            in1 => \N__17571\,
            in2 => \_gnd_net_\,
            in3 => \N__17679\,
            lcout => \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_rx_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10702\,
            in1 => \N__10132\,
            in2 => \_gnd_net_\,
            in3 => \N__10117\,
            lcout => \spi_slave_1.bitcnt_rxZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \spi_slave_1.bitcnt_rx_cry_0\,
            clk => \N__27448\,
            ce => \N__12064\,
            sr => \N__27100\
        );

    \spi_slave_1.bitcnt_rx_1_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10710\,
            in1 => \N__10114\,
            in2 => \_gnd_net_\,
            in3 => \N__10102\,
            lcout => \spi_slave_1.bitcnt_rxZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_slave_1.bitcnt_rx_cry_0\,
            carryout => \spi_slave_1.bitcnt_rx_cry_1\,
            clk => \N__27448\,
            ce => \N__12064\,
            sr => \N__27100\
        );

    \spi_slave_1.bitcnt_rx_2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10703\,
            in1 => \N__10099\,
            in2 => \_gnd_net_\,
            in3 => \N__10087\,
            lcout => \spi_slave_1.bitcnt_rxZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_slave_1.bitcnt_rx_cry_1\,
            carryout => \spi_slave_1.bitcnt_rx_cry_2\,
            clk => \N__27448\,
            ce => \N__12064\,
            sr => \N__27100\
        );

    \spi_slave_1.bitcnt_rx_3_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10711\,
            in1 => \N__10192\,
            in2 => \_gnd_net_\,
            in3 => \N__10180\,
            lcout => \spi_slave_1.bitcnt_rxZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_1.bitcnt_rx_cry_2\,
            carryout => \spi_slave_1.bitcnt_rx_cry_3\,
            clk => \N__27448\,
            ce => \N__12064\,
            sr => \N__27100\
        );

    \spi_slave_1.bitcnt_rx_4_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10704\,
            in1 => \N__10174\,
            in2 => \_gnd_net_\,
            in3 => \N__10177\,
            lcout => \spi_slave_1.bitcnt_rxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27448\,
            ce => \N__12064\,
            sr => \N__27100\
        );

    \spi_slave_1.miso_en_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__10159\,
            in1 => \N__10885\,
            in2 => \N__11877\,
            in3 => \N__10861\,
            lcout => miso_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27454\,
            ce => 'H',
            sr => \N__27110\
        );

    \sb_translator_1.instr_tmp_17_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__11335\,
            in1 => \N__22075\,
            in2 => \N__14667\,
            in3 => \N__16852\,
            lcout => \sb_translator_1.instr_tmpZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27454\,
            ce => 'H',
            sr => \N__27110\
        );

    \spi_slave_1.un1_bitcnt_tx_1_cry_0_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18512\,
            in2 => \N__10783\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \spi_slave_1.un1_bitcnt_tx_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_LUT4_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11941\,
            in2 => \_gnd_net_\,
            in3 => \N__10153\,
            lcout => \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_1.un1_bitcnt_tx_1_cry_0\,
            carryout => \spi_slave_1.un1_bitcnt_tx_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_LUT4_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11694\,
            in2 => \_gnd_net_\,
            in3 => \N__10150\,
            lcout => \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_1.un1_bitcnt_tx_1_cry_1\,
            carryout => \spi_slave_1.un1_bitcnt_tx_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_3_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27159\,
            in1 => \N__10860\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => \spi_slave_1.bitcnt_txZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_1.un1_bitcnt_tx_1_cry_2\,
            carryout => \spi_slave_1.un1_bitcnt_tx_1_cry_3\,
            clk => \N__27464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110111010"
        )
    port map (
            in0 => \N__27158\,
            in1 => \N__10914\,
            in2 => \N__18580\,
            in3 => \N__10144\,
            lcout => \spi_slave_1.bitcnt_txZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001110"
        )
    port map (
            in0 => \N__11695\,
            in1 => \N__27157\,
            in2 => \N__10921\,
            in3 => \N__10204\,
            lcout => \spi_slave_1.bitcnt_txZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_1_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111110010"
        )
    port map (
            in0 => \N__11942\,
            in1 => \N__10915\,
            in2 => \N__27160\,
            in3 => \N__10198\,
            lcout => \spi_slave_1.bitcnt_txZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.mosi_data_in_18_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12087\,
            in1 => \N__12186\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_19_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12324\,
            in1 => \_gnd_net_\,
            in2 => \N__12224\,
            in3 => \N__10263\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_20_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10251\,
            in1 => \N__12190\,
            in2 => \_gnd_net_\,
            in3 => \N__12325\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_21_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12326\,
            in1 => \_gnd_net_\,
            in2 => \N__12225\,
            in3 => \N__10239\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_22_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10227\,
            in1 => \N__12194\,
            in2 => \_gnd_net_\,
            in3 => \N__12327\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_23_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12328\,
            in1 => \_gnd_net_\,
            in2 => \N__12226\,
            in3 => \N__10215\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_8_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13198\,
            in1 => \N__12198\,
            in2 => \_gnd_net_\,
            in3 => \N__12329\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_in_9_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12330\,
            in1 => \_gnd_net_\,
            in2 => \N__12227\,
            in3 => \N__12015\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27421\,
            ce => \N__12062\,
            sr => \N__27065\
        );

    \spi_slave_1.mosi_data_out_17_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12088\,
            lcout => mosi_data_out_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_23_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10270\,
            lcout => mosi_data_out_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_18_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10264\,
            lcout => mosi_data_out_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_19_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10252\,
            lcout => mosi_data_out_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_1_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => mosi_data_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_20_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10240\,
            lcout => mosi_data_out_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_21_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10228\,
            lcout => mosi_data_out_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \spi_slave_1.mosi_data_out_22_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10216\,
            lcout => mosi_data_out_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27422\,
            ce => \N__18424\,
            sr => \N__27067\
        );

    \sb_translator_1.cnt_10_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__22763\,
            in1 => \N__17094\,
            in2 => \N__17220\,
            in3 => \N__10330\,
            lcout => \sb_translator_1.cntZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_2_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17090\,
            in1 => \N__17177\,
            in2 => \N__22786\,
            in3 => \N__10324\,
            lcout => \sb_translator_1.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_3_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__22764\,
            in1 => \N__17095\,
            in2 => \N__17221\,
            in3 => \N__10318\,
            lcout => \sb_translator_1.cntZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17091\,
            in1 => \N__17178\,
            in2 => \N__22787\,
            in3 => \N__10312\,
            lcout => \sb_translator_1.cntZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_5_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__22765\,
            in1 => \N__17096\,
            in2 => \N__17222\,
            in3 => \N__10306\,
            lcout => \sb_translator_1.cntZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_6_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17092\,
            in1 => \N__17179\,
            in2 => \N__22788\,
            in3 => \N__10300\,
            lcout => \sb_translator_1.cntZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_7_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__22766\,
            in1 => \N__17097\,
            in2 => \N__17223\,
            in3 => \N__10294\,
            lcout => \sb_translator_1.cntZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.cnt_8_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17093\,
            in1 => \N__17180\,
            in2 => \N__22789\,
            in3 => \N__10288\,
            lcout => \sb_translator_1.cntZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27427\,
            ce => 'H',
            sr => \N__27070\
        );

    \sb_translator_1.state_5_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17199\,
            in1 => \N__22735\,
            in2 => \_gnd_net_\,
            in3 => \N__17104\,
            lcout => \sb_translator_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_RNO_0_0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12512\,
            in2 => \_gnd_net_\,
            in3 => \N__16881\,
            lcout => OPEN,
            ltout => \sb_translator_1.cnt_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001000011110000"
        )
    port map (
            in0 => \N__17196\,
            in1 => \N__22734\,
            in2 => \N__10432\,
            in3 => \N__17103\,
            lcout => \sb_translator_1.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_13_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17098\,
            in1 => \N__17200\,
            in2 => \N__22779\,
            in3 => \N__10429\,
            lcout => \sb_translator_1.cntZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_14_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__17197\,
            in1 => \N__17101\,
            in2 => \N__22782\,
            in3 => \N__10408\,
            lcout => \sb_translator_1.cntZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_15_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17099\,
            in1 => \N__17201\,
            in2 => \N__22780\,
            in3 => \N__10387\,
            lcout => \sb_translator_1.cntZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_16_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__17198\,
            in1 => \N__17102\,
            in2 => \N__22783\,
            in3 => \N__10366\,
            lcout => \sb_translator_1.cntZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_1_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17100\,
            in1 => \N__17202\,
            in2 => \N__22781\,
            in3 => \N__10348\,
            lcout => \sb_translator_1.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27429\,
            ce => 'H',
            sr => \N__27074\
        );

    \sb_translator_1.cnt_11_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17105\,
            in1 => \N__22760\,
            in2 => \N__17227\,
            in3 => \N__10342\,
            lcout => \sb_translator_1.cntZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27435\,
            ce => 'H',
            sr => \N__27077\
        );

    \sb_translator_1.cnt_12_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011011100000000"
        )
    port map (
            in0 => \N__22759\,
            in1 => \N__17107\,
            in2 => \N__17234\,
            in3 => \N__10336\,
            lcout => \sb_translator_1.cntZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27435\,
            ce => 'H',
            sr => \N__27077\
        );

    \sb_translator_1.cnt_9_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011100000000"
        )
    port map (
            in0 => \N__17106\,
            in1 => \N__22761\,
            in2 => \N__17228\,
            in3 => \N__10570\,
            lcout => \sb_translator_1.cntZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27435\,
            ce => 'H',
            sr => \N__27077\
        );

    \sb_translator_1.cnt_RNIJ7EF_1_9_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__22057\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__10557\,
            lcout => \sb_translator_1.cnt_RNIJ7EF_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIJ7EF_2_9_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__10558\,
            in1 => \_gnd_net_\,
            in2 => \N__10529\,
            in3 => \N__22059\,
            lcout => \sb_translator_1.cnt_RNIJ7EF_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIJ7EF_0_9_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22058\,
            in1 => \N__10522\,
            in2 => \_gnd_net_\,
            in3 => \N__10559\,
            lcout => \sb_translator_1.N_1088\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNIJ7EF_9_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__10560\,
            in1 => \_gnd_net_\,
            in2 => \N__10530\,
            in3 => \N__22060\,
            lcout => \sb_translator_1.N_1092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_tmp_22_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__22061\,
            in1 => \N__17203\,
            in2 => \N__10630\,
            in3 => \N__16864\,
            lcout => \sb_translator_1.instr_tmpZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27435\,
            ce => 'H',
            sr => \N__27077\
        );

    \sb_translator_1.instr_out_18_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10491\,
            lcout => miso_data_in_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_19_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10476\,
            lcout => miso_data_in_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_20_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => miso_data_in_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_21_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10446\,
            lcout => miso_data_in_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_22_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10629\,
            lcout => miso_data_in_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_23_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10614\,
            lcout => miso_data_in_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_8_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15621\,
            lcout => miso_data_in_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \sb_translator_1.instr_out_9_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => miso_data_in_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27441\,
            ce => \N__23993\,
            sr => \N__27082\
        );

    \spi_slave_1.miso_data_out_19_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.miso_data_outZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_20_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10594\,
            lcout => \spi_slave_1.miso_data_outZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_21_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10588\,
            lcout => \spi_slave_1.miso_data_outZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_22_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10582\,
            lcout => \spi_slave_1.miso_data_outZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_23_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10576\,
            lcout => \spi_slave_1.miso_data_outZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_5_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24277\,
            lcout => \spi_slave_1.miso_data_outZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_8_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10717\,
            lcout => \spi_slave_1.miso_data_outZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_4_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24013\,
            lcout => \spi_slave_1.miso_data_outZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27449\,
            ce => \N__14547\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.clk_RNIDBLL_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12146\,
            lcout => \spi_slave_1.clk_pos_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_18_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__11524\,
            in1 => \N__18582\,
            in2 => \N__10687\,
            in3 => \N__18504\,
            lcout => OPEN,
            ltout => \spi_slave_1.m81_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_16_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__18506\,
            in1 => \N__10678\,
            in2 => \N__10672\,
            in3 => \N__10669\,
            lcout => \spi_slave_1.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_15_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__10663\,
            in1 => \N__18583\,
            in2 => \N__10657\,
            in3 => \N__18505\,
            lcout => OPEN,
            ltout => \spi_slave_1.m60_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_10_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__18507\,
            in1 => \N__10648\,
            in2 => \N__10642\,
            in3 => \N__11770\,
            lcout => \spi_slave_1.miso_RNOZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.clk_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.clkZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.clk_RNIFQ8K3_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__12111\,
            in1 => \N__12267\,
            in2 => \N__11864\,
            in3 => \N__10830\,
            lcout => \spi_slave_1.bitcnt_tx10\,
            ltout => \spi_slave_1.bitcnt_tx10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_0_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011110"
        )
    port map (
            in0 => \N__18510\,
            in1 => \N__27153\,
            in2 => \N__10774\,
            in3 => \N__10919\,
            lcout => \spi_slave_1.bitcnt_txZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_2_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12112\,
            in1 => \N__12268\,
            in2 => \_gnd_net_\,
            in3 => \N__10831\,
            lcout => \spi_slave_1.N_96_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_7_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__18509\,
            in1 => \N__10771\,
            in2 => \_gnd_net_\,
            in3 => \N__11758\,
            lcout => \spi_slave_1.miso_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.clk_1_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12269\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.clkZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_RNIQORT2_3_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10883\,
            in1 => \N__10762\,
            in2 => \N__11863\,
            in3 => \N__10859\,
            lcout => \spi_slave_1.miso_data_out_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_17_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101000100"
        )
    port map (
            in0 => \N__11512\,
            in1 => \N__18508\,
            in2 => \N__14566\,
            in3 => \N__11722\,
            lcout => \spi_slave_1.miso_RNOZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_11_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__11934\,
            in1 => \N__10744\,
            in2 => \N__11697\,
            in3 => \N__10735\,
            lcout => OPEN,
            ltout => \spi_slave_1.m48_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__18454\,
            in1 => \N__10729\,
            in2 => \N__10720\,
            in3 => \N__11935\,
            lcout => OPEN,
            ltout => \spi_slave_1.N_49_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__10863\,
            in1 => \_gnd_net_\,
            in2 => \N__10939\,
            in3 => \N__11896\,
            lcout => OPEN,
            ltout => \spi_slave_1.N_25_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__11841\,
            in1 => \_gnd_net_\,
            in2 => \N__10936\,
            in3 => \N__10933\,
            lcout => \spi_slave_1.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_RNIP9N23_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11274\,
            in2 => \_gnd_net_\,
            in3 => \N__10920\,
            lcout => \spi_slave_1.bitcnt_tx_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_0_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000101111"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__10864\,
            in2 => \N__11862\,
            in3 => \N__10891\,
            lcout => \spi_slave_1.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_RNIJITN1_2_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11933\,
            in1 => \N__18563\,
            in2 => \N__11696\,
            in3 => \N__18511\,
            lcout => \spi_slave_1.N_94_mux\,
            ltout => \spi_slave_1.N_94_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.bitcnt_tx_RNIGFSJ2_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__18564\,
            in1 => \_gnd_net_\,
            in2 => \N__10867\,
            in3 => \N__10862\,
            lcout => \spi_slave_1.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__10806\,
            in1 => \N__10822\,
            in2 => \_gnd_net_\,
            in3 => \N__10816\,
            lcout => miso,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27480\,
            ce => 'H',
            sr => \N__27113\
        );

    \spi_slave_1.clk_RNIVAC01_1_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__12202\,
            in1 => \N__11878\,
            in2 => \_gnd_net_\,
            in3 => \N__12348\,
            lcout => \spi_slave_1.bitcnt_rxe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_6_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.num_ledsZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27425\,
            ce => \N__22362\,
            sr => \N__27063\
        );

    \sb_translator_1.num_leds_5_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13855\,
            lcout => \sb_translator_1.num_ledsZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27425\,
            ce => \N__22362\,
            sr => \N__27063\
        );

    \sb_translator_1.num_leds_RNIN668_0_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19104\,
            in2 => \N__19042\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.un1_num_leds_n_1\,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_1_c_RNIDRFK_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19041\,
            in2 => \N__19071\,
            in3 => \N__11023\,
            lcout => \sb_translator_1.un1_num_leds_n_2\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_1\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_2_c_RNIGVGK_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19061\,
            in2 => \N__18685\,
            in3 => \N__11008\,
            lcout => \sb_translator_1.un1_num_leds_n_3\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_2\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_3_c_RNIJ3IK_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18680\,
            in2 => \N__18643\,
            in3 => \N__10996\,
            lcout => \sb_translator_1.un1_num_leds_n_4\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_3\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_4_c_RNIM7JK_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18634\,
            in2 => \N__18402\,
            in3 => \N__10984\,
            lcout => \sb_translator_1.un1_num_leds_n_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_4\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_5_c_RNIPBKK_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18392\,
            in2 => \N__18795\,
            in3 => \N__10969\,
            lcout => \sb_translator_1.un1_num_leds_n_6\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_5\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_6_c_RNISFLK_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18785\,
            in2 => \N__18753\,
            in3 => \N__10957\,
            lcout => \sb_translator_1.un1_num_leds_n_7\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_6\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_7_c_RNIVJMK_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18749\,
            in2 => \N__18728\,
            in3 => \N__10942\,
            lcout => \sb_translator_1.un1_num_leds_n_8\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_7\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_8_c_RNI2ONK_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18722\,
            in2 => \N__15934\,
            in3 => \N__11134\,
            lcout => \sb_translator_1.un1_num_leds_n_9\,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_9_c_RNIC3RN_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15932\,
            in2 => \N__15874\,
            in3 => \N__11122\,
            lcout => \sb_translator_1.un1_num_leds_n_10\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_9\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_10_c_RNITFLI_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15872\,
            in2 => \N__15901\,
            in3 => \N__11107\,
            lcout => \sb_translator_1.un1_num_leds_n_11\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_10\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_11_c_RNI0KMI_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15900\,
            in2 => \N__20876\,
            in3 => \N__11095\,
            lcout => \sb_translator_1.un1_num_leds_n_12\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_11\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_12_c_RNI3ONI_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20870\,
            in2 => \N__20775\,
            in3 => \N__11083\,
            lcout => \sb_translator_1.un1_num_leds_n_13\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_12\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_13_c_RNI6SOI_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20765\,
            in2 => \N__20802\,
            in3 => \N__11071\,
            lcout => \sb_translator_1.un1_num_leds_n_14\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_13\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_14_c_RNI90QI_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20798\,
            in2 => \N__20962\,
            in3 => \N__11059\,
            lcout => \sb_translator_1.un1_num_leds_n_15\,
            ltout => OPEN,
            carryin => \sb_translator_1.un1_num_leds_0_cry_14\,
            carryout => \sb_translator_1.un1_num_leds_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.un1_num_leds_0_cry_15_c_RNIQ9LB_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20961\,
            in2 => \_gnd_net_\,
            in3 => \N__11056\,
            lcout => \sb_translator_1.un1_num_leds_n_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.mosi_data_in_0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11887\,
            in1 => \N__12228\,
            in2 => \_gnd_net_\,
            in3 => \N__12357\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_1_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12358\,
            in1 => \_gnd_net_\,
            in2 => \N__12244\,
            in3 => \N__13167\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_2_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11154\,
            in1 => \N__12232\,
            in2 => \_gnd_net_\,
            in3 => \N__12359\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_3_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12360\,
            in1 => \_gnd_net_\,
            in2 => \N__12245\,
            in3 => \N__12375\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_4_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12387\,
            in1 => \N__12236\,
            in2 => \_gnd_net_\,
            in3 => \N__12361\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_5_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12362\,
            in1 => \_gnd_net_\,
            in2 => \N__12246\,
            in3 => \N__13179\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_6_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13221\,
            in1 => \N__12240\,
            in2 => \_gnd_net_\,
            in3 => \N__12363\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \spi_slave_1.mosi_data_in_7_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12364\,
            in1 => \_gnd_net_\,
            in2 => \N__12247\,
            in3 => \N__13209\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27436\,
            ce => \N__12063\,
            sr => \N__27071\
        );

    \sb_translator_1.instr_tmp_5_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22043\,
            in1 => \N__13848\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.instr_tmpZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27444\,
            ce => \N__16971\,
            sr => \N__27075\
        );

    \sb_translator_1.instr_tmp_6_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22042\,
            in2 => \_gnd_net_\,
            in3 => \N__13689\,
            lcout => \sb_translator_1.instr_tmpZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27444\,
            ce => \N__16971\,
            sr => \N__27075\
        );

    \sb_translator_1.instr_tmp_7_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22044\,
            in1 => \N__13509\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.instr_tmpZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27444\,
            ce => \N__16971\,
            sr => \N__27075\
        );

    \reset_n_input_RNIVGR4_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11281\,
            lcout => reset_n_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_3_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__13920\,
            in1 => \N__13947\,
            in2 => \N__17536\,
            in3 => \N__13301\,
            lcout => ram_we_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.ram_we_13_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17761\,
            in1 => \N__14048\,
            in2 => \N__11376\,
            in3 => \N__13919\,
            lcout => ram_we_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.cnt_RNILAHE_0_10_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__17359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17311\,
            lcout => \sb_translator_1.cnt_RNILAHE_0Z0Z_10\,
            ltout => \sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_5_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__13945\,
            in1 => \N__17794\,
            in2 => \N__11200\,
            in3 => \N__13921\,
            lcout => ram_we_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.ram_we_7_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13922\,
            in1 => \N__13946\,
            in2 => \N__17275\,
            in3 => \N__16950\,
            lcout => ram_we_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.ram_we_9_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16108\,
            in1 => \N__14283\,
            in2 => \N__11377\,
            in3 => \N__13923\,
            lcout => ram_we_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.cnt_RNILAHE_1_10_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17312\,
            lcout => \sb_translator_1.cnt_RNILAHE_1Z0Z_10\,
            ltout => \sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_11_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__11369\,
            in1 => \N__16915\,
            in2 => \N__11356\,
            in3 => \N__13918\,
            lcout => ram_we_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27450\,
            ce => \N__16785\,
            sr => \N__27078\
        );

    \sb_translator_1.state_RNIHS98_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22049\,
            lcout => \sb_translator_1.state_RNIHS98Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNIHS98_0_0_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__22048\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11328\,
            lcout => \sb_translator_1.state_RNIHS98_0Z0Z_0\,
            ltout => \sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_6_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__15841\,
            in1 => \N__21313\,
            in2 => \N__11338\,
            in3 => \N__16951\,
            lcout => ram_sel_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27457\,
            ce => \N__17482\,
            sr => \N__27083\
        );

    \sb_translator_1.state_RNIQIHP_0_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__22045\,
            in1 => \N__16860\,
            in2 => \_gnd_net_\,
            in3 => \N__22417\,
            lcout => \sb_translator_1.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNO_0_0_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16862\,
            in1 => \N__22602\,
            in2 => \_gnd_net_\,
            in3 => \N__22046\,
            lcout => \sb_translator_1.N_729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNI9ILJ_0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17232\,
            in1 => \N__22053\,
            in2 => \N__22603\,
            in3 => \N__11331\,
            lcout => \sb_translator_1.state_RNI9ILJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNI9ILJ_0_0_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11330\,
            in1 => \N__22598\,
            in2 => \N__22074\,
            in3 => \N__17233\,
            lcout => \sb_translator_1.state_RNI9ILJ_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNII30C_0_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__22047\,
            in1 => \_gnd_net_\,
            in2 => \N__17236\,
            in3 => \N__16861\,
            lcout => \sb_translator_1.state_RNII30CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_a3_2_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11299\,
            lcout => OPEN,
            ltout => \demux.N_877_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_9_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14485\,
            in1 => \N__11503\,
            in2 => \N__11494\,
            in3 => \N__11476\,
            lcout => \demux.N_418_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_6_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__19645\,
            in1 => \N__11491\,
            in2 => \N__24360\,
            in3 => \N__11482\,
            lcout => \demux.N_418_i_0_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_a3_2_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11470\,
            in2 => \_gnd_net_\,
            in3 => \N__17946\,
            lcout => OPEN,
            ltout => \demux.N_835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_9_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__11452\,
            in1 => \N__14484\,
            in2 => \N__11446\,
            in3 => \N__11425\,
            lcout => \demux.N_421_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_6_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__11443\,
            in1 => \N__24349\,
            in2 => \N__11437\,
            in3 => \N__19643\,
            lcout => \demux.N_421_i_0_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_a3_1_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19644\,
            in1 => \N__11419\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \demux.N_890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_a3_1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11413\,
            in2 => \_gnd_net_\,
            in3 => \N__19642\,
            lcout => \demux.N_423_i_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_6_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__17944\,
            in1 => \N__11407\,
            in2 => \N__21069\,
            in3 => \N__11389\,
            lcout => OPEN,
            ltout => \demux.N_417_i_0_o2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_9_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__11662\,
            in1 => \N__14471\,
            in2 => \N__11650\,
            in3 => \N__11647\,
            lcout => \demux.N_417_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_a3_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11641\,
            in2 => \_gnd_net_\,
            in3 => \N__19653\,
            lcout => \demux.N_419_i_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_6_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__11635\,
            in1 => \N__17943\,
            in2 => \N__11623\,
            in3 => \N__21052\,
            lcout => OPEN,
            ltout => \demux.N_419_i_0_o2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_9_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14470\,
            in1 => \N__11602\,
            in2 => \N__11587\,
            in3 => \N__11584\,
            lcout => \demux.N_419_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_a3_1_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11578\,
            lcout => \demux.N_420_i_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_6_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__17945\,
            in1 => \N__11572\,
            in2 => \N__21070\,
            in3 => \N__11554\,
            lcout => OPEN,
            ltout => \demux.N_420_i_0_o2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_9_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__11542\,
            in1 => \N__14472\,
            in2 => \N__11533\,
            in3 => \N__11530\,
            lcout => \demux.N_420_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_6_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23533\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.miso_data_outZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24022\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.miso_data_outZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_3_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.miso_data_outZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_7_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23671\,
            lcout => \spi_slave_1.miso_data_outZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_18_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11749\,
            lcout => \spi_slave_1.miso_data_outZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_2_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17248\,
            lcout => \spi_slave_1.miso_data_outZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27481\,
            ce => \N__14546\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_19_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__11737\,
            in1 => \N__18571\,
            in2 => \N__11731\,
            in3 => \N__18521\,
            lcout => \spi_slave_1.m72_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_14_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_1.miso_data_outZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27489\,
            ce => \N__14539\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_13_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14698\,
            lcout => \spi_slave_1.miso_data_outZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27489\,
            ce => \N__14539\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_12_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__18522\,
            in1 => \N__11710\,
            in2 => \_gnd_net_\,
            in3 => \N__11704\,
            lcout => OPEN,
            ltout => \spi_slave_1.miso_RNOZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_8_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__11698\,
            in1 => \N__11943\,
            in2 => \N__11665\,
            in3 => \N__17962\,
            lcout => OPEN,
            ltout => \spi_slave_1.m27_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_4_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__11944\,
            in1 => \N__18604\,
            in2 => \N__11911\,
            in3 => \N__11908\,
            lcout => \spi_slave_1.N_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.mosi_buffer_1_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11869\,
            in2 => \_gnd_net_\,
            in3 => \N__11776\,
            lcout => \spi_slave_1.mosi_bufferZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27494\,
            ce => 'H',
            sr => \N__27114\
        );

    \spi_slave_1.mosi_buffer_0_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11791\,
            lcout => \spi_slave_1.mosi_bufferZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27494\,
            ce => 'H',
            sr => \N__27114\
        );

    \spi_slave_1.mosi_data_in_10_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__12170\,
            in2 => \_gnd_net_\,
            in3 => \N__12349\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_11_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12350\,
            in1 => \_gnd_net_\,
            in2 => \N__12220\,
            in3 => \N__12003\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_12_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11991\,
            in1 => \N__12174\,
            in2 => \_gnd_net_\,
            in3 => \N__12351\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_13_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12352\,
            in1 => \_gnd_net_\,
            in2 => \N__12221\,
            in3 => \N__11979\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_14_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11967\,
            in1 => \N__12178\,
            in2 => \_gnd_net_\,
            in3 => \N__12353\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_15_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12354\,
            in1 => \_gnd_net_\,
            in2 => \N__12222\,
            in3 => \N__11955\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_16_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18438\,
            in1 => \N__12182\,
            in2 => \_gnd_net_\,
            in3 => \N__12355\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_in_17_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12356\,
            in1 => \_gnd_net_\,
            in2 => \N__12223\,
            in3 => \N__12399\,
            lcout => \spi_slave_1.mosi_data_inZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27426\,
            ce => \N__12061\,
            sr => \N__27064\
        );

    \spi_slave_1.mosi_data_out_9_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12046\,
            lcout => mosi_data_out_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_8_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12022\,
            lcout => mosi_data_out_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_10_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12004\,
            lcout => mosi_data_out_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_11_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11992\,
            lcout => mosi_data_out_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_12_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11980\,
            lcout => mosi_data_out_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_13_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11968\,
            lcout => mosi_data_out_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \spi_slave_1.mosi_data_out_14_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11956\,
            lcout => mosi_data_out_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27428\,
            ce => \N__18426\,
            sr => \N__27066\
        );

    \sb_translator_1.num_leds_11_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14644\,
            lcout => \sb_translator_1.num_ledsZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_12_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22578\,
            lcout => \sb_translator_1.num_ledsZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_13_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14605\,
            lcout => \sb_translator_1.num_ledsZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_14_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22521\,
            lcout => \sb_translator_1.num_ledsZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_2_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15961\,
            lcout => \sb_translator_1.num_ledsZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_3_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17029\,
            lcout => \sb_translator_1.num_ledsZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_4_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17002\,
            lcout => \sb_translator_1.num_ledsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_7_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13513\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.num_ledsZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27432\,
            ce => \N__22349\,
            sr => \N__27068\
        );

    \sb_translator_1.num_leds_RNITOUT_8_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \N__20476\,
            in1 => \N__21356\,
            in2 => \N__15933\,
            in3 => \N__18717\,
            lcout => \sb_translator_1.num_leds_RNITOUTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNI0EVE_8_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__18718\,
            in1 => \_gnd_net_\,
            in2 => \N__21364\,
            in3 => \N__15928\,
            lcout => \sb_translator_1.num_leds_RNI0EVEZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_8_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.num_ledsZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27437\,
            ce => \N__22363\,
            sr => \N__27072\
        );

    \sb_translator_1.num_leds_9_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12484\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.num_ledsZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27437\,
            ce => \N__22363\,
            sr => \N__27072\
        );

    \sb_translator_1.addr_out_RNO_0_0_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12531\,
            in1 => \N__22997\,
            in2 => \_gnd_net_\,
            in3 => \N__12517\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_RNO_0_1_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22998\,
            in1 => \N__12483\,
            in2 => \_gnd_net_\,
            in3 => \N__12472\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_RNO_0_2_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12414\,
            in1 => \N__22999\,
            in2 => \_gnd_net_\,
            in3 => \N__12442\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_10_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12415\,
            lcout => \sb_translator_1.num_ledsZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27437\,
            ce => \N__22363\,
            sr => \N__27072\
        );

    \spi_slave_1.mosi_data_out_16_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12403\,
            lcout => mosi_data_out_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_3_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12388\,
            lcout => mosi_data_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12376\,
            lcout => mosi_data_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_5_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13222\,
            lcout => mosi_data_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_6_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13210\,
            lcout => mosi_data_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_7_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13194\,
            lcout => mosi_data_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_4_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13180\,
            lcout => mosi_data_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \spi_slave_1.mosi_data_out_0_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13168\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => mosi_data_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27445\,
            ce => \N__18425\,
            sr => \N__27076\
        );

    \sb_translator_1.data_out_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16022\,
            in1 => \N__21993\,
            in2 => \_gnd_net_\,
            in3 => \N__16003\,
            lcout => ram_data_in_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21989\,
            in1 => \N__15967\,
            in2 => \_gnd_net_\,
            in3 => \N__15989\,
            lcout => ram_data_in_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_2_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15940\,
            in1 => \N__15956\,
            in2 => \_gnd_net_\,
            in3 => \N__21994\,
            lcout => ram_data_in_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21990\,
            in1 => \N__17008\,
            in2 => \_gnd_net_\,
            in3 => \N__17024\,
            lcout => ram_data_in_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17000\,
            in1 => \N__21995\,
            in2 => \_gnd_net_\,
            in3 => \N__16981\,
            lcout => ram_data_in_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_5_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21991\,
            in1 => \N__13861\,
            in2 => \_gnd_net_\,
            in3 => \N__13847\,
            lcout => ram_data_in_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13702\,
            in1 => \N__13688\,
            in2 => \_gnd_net_\,
            in3 => \N__21996\,
            lcout => ram_data_in_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.data_out_7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21992\,
            in1 => \N__13519\,
            in2 => \_gnd_net_\,
            in3 => \N__13508\,
            lcout => ram_data_in_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27451\,
            ce => \N__16789\,
            sr => \N__27079\
        );

    \sb_translator_1.ram_we_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__14011\,
            in1 => \N__16099\,
            in2 => \N__17728\,
            in3 => \N__13990\,
            lcout => ram_we_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13987\,
            in1 => \N__17529\,
            in2 => \N__13306\,
            in3 => \N__14014\,
            lcout => ram_we_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_10_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__13302\,
            in2 => \N__16918\,
            in3 => \N__13991\,
            lcout => ram_we_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_8_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__13989\,
            in1 => \N__13254\,
            in2 => \N__16104\,
            in3 => \N__14282\,
            lcout => ram_we_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_12_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17757\,
            in1 => \N__14049\,
            in2 => \N__13255\,
            in3 => \N__13992\,
            lcout => ram_we_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13988\,
            in1 => \N__17792\,
            in2 => \N__14053\,
            in3 => \N__14012\,
            lcout => ram_we_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14013\,
            in1 => \N__16945\,
            in2 => \N__17265\,
            in3 => \N__13993\,
            lcout => ram_we_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_we_1_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17727\,
            in1 => \N__13951\,
            in2 => \N__16103\,
            in3 => \N__13924\,
            lcout => ram_we_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27458\,
            ce => \N__16784\,
            sr => \N__27084\
        );

    \sb_translator_1.ram_sel_11_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16071\,
            in1 => \N__16916\,
            in2 => \N__13873\,
            in3 => \N__14343\,
            lcout => ram_sel_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27466\,
            ce => \N__17483\,
            sr => \N__27089\
        );

    \sb_translator_1.cnt_leds_RNI1VFQ_9_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__21362\,
            in1 => \_gnd_net_\,
            in2 => \N__21418\,
            in3 => \N__22052\,
            lcout => \sb_translator_1.N_1091\,
            ltout => \sb_translator_1.N_1091_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_13_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17750\,
            in1 => \N__15809\,
            in2 => \N__13879\,
            in3 => \N__14344\,
            lcout => ram_sel_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27466\,
            ce => \N__17483\,
            sr => \N__27089\
        );

    \sb_translator_1.cnt_leds_RNI1VFQ_0_9_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__21361\,
            in1 => \_gnd_net_\,
            in2 => \N__21417\,
            in3 => \N__22051\,
            lcout => \sb_translator_1.N_1089\,
            ltout => \sb_translator_1.N_1089_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_10_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16070\,
            in1 => \N__14295\,
            in2 => \N__13876\,
            in3 => \N__16917\,
            lcout => ram_sel_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27466\,
            ce => \N__17483\,
            sr => \N__27089\
        );

    \sb_translator_1.ram_sel_9_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14342\,
            in1 => \N__16038\,
            in2 => \N__14281\,
            in3 => \N__13872\,
            lcout => ram_sel_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27466\,
            ce => \N__17483\,
            sr => \N__27089\
        );

    \sb_translator_1.cnt_leds_RNI1VFQ_1_9_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__22050\,
            in1 => \N__21409\,
            in2 => \_gnd_net_\,
            in3 => \N__21360\,
            lcout => \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9\,
            ltout => \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_7_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__14341\,
            in1 => \N__16946\,
            in2 => \N__14218\,
            in3 => \N__15840\,
            lcout => ram_sel_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27466\,
            ce => \N__17483\,
            sr => \N__27089\
        );

    \demux.N_422_i_0_o2_6_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__14215\,
            in1 => \N__21060\,
            in2 => \N__14200\,
            in3 => \N__17936\,
            lcout => OPEN,
            ltout => \demux.N_422_i_0_o2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_9_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14182\,
            in1 => \N__14477\,
            in2 => \N__14170\,
            in3 => \N__14104\,
            lcout => \demux.N_422_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_6_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__14167\,
            in1 => \N__21059\,
            in2 => \N__14152\,
            in3 => \N__17935\,
            lcout => OPEN,
            ltout => \demux.N_423_i_0_o2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_9_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14137\,
            in1 => \N__14476\,
            in2 => \N__14125\,
            in3 => \N__14122\,
            lcout => \demux.N_423_i_0_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_a3_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14116\,
            in2 => \_gnd_net_\,
            in3 => \N__19651\,
            lcout => \demux.N_422_i_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_6_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__17937\,
            in1 => \N__14098\,
            in2 => \N__21071\,
            in3 => \N__14083\,
            lcout => OPEN,
            ltout => \demux.N_424_i_0_o2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_9_0_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14478\,
            in1 => \N__14071\,
            in2 => \N__14056\,
            in3 => \N__14371\,
            lcout => \demux.N_424_i_0_o2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a3_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14383\,
            lcout => \demux.N_424_i_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__21310\,
            in1 => \N__17719\,
            in2 => \N__16054\,
            in3 => \N__14310\,
            lcout => ram_sel_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_2_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14312\,
            in1 => \N__21312\,
            in2 => \N__17527\,
            in3 => \N__16077\,
            lcout => ram_sel_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14364\,
            in1 => \N__14346\,
            in2 => \N__16053\,
            in3 => \N__17720\,
            lcout => ram_sel_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_3_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14345\,
            in1 => \N__14365\,
            in2 => \N__17528\,
            in3 => \N__16078\,
            lcout => ram_sel_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_5_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__14363\,
            in1 => \N__17788\,
            in2 => \N__14350\,
            in3 => \N__15819\,
            lcout => ram_sel_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_4_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14313\,
            in1 => \N__21311\,
            in2 => \N__17793\,
            in3 => \N__15820\,
            lcout => ram_sel_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_12_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__17749\,
            in1 => \N__15818\,
            in2 => \N__14233\,
            in3 => \N__14311\,
            lcout => ram_sel_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \sb_translator_1.ram_sel_8_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__14314\,
            in1 => \N__16049\,
            in2 => \N__14284\,
            in3 => \N__14232\,
            lcout => ram_sel_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27482\,
            ce => \N__17494\,
            sr => \N__27101\
        );

    \demux.N_424_i_0_o2_11_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17854\,
            in2 => \_gnd_net_\,
            in3 => \N__17875\,
            lcout => \demux.N_236\,
            ltout => \demux.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_16_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14436\,
            in2 => \N__14491\,
            in3 => \N__14415\,
            lcout => \demux.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_14_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19806\,
            in2 => \_gnd_net_\,
            in3 => \N__19752\,
            lcout => \demux.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_10_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14437\,
            in2 => \_gnd_net_\,
            in3 => \N__14416\,
            lcout => \demux.N_235\,
            ltout => \demux.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17857\,
            in1 => \N__17879\,
            in2 => \N__14488\,
            in3 => \N__17891\,
            lcout => \demux.N_424_i_0_a2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_6_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__17893\,
            in1 => \N__14442\,
            in2 => \N__19602\,
            in3 => \N__14419\,
            lcout => \demux.N_424_i_0_a2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14418\,
            in1 => \N__19595\,
            in2 => \N__14443\,
            in3 => \N__17892\,
            lcout => \demux.N_424_i_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__17855\,
            in1 => \N__14438\,
            in2 => \N__17881\,
            in3 => \N__14417\,
            lcout => \demux.N_424_i_0_o2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17806\,
            lcout => \spi_slave_1.miso_data_outZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_9_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14398\,
            lcout => \spi_slave_1.miso_data_outZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_10_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14509\,
            lcout => \spi_slave_1.miso_data_outZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_11_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14503\,
            lcout => \spi_slave_1.miso_data_outZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_12_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14497\,
            lcout => \spi_slave_1.miso_data_outZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_15_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14686\,
            lcout => \spi_slave_1.miso_data_outZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_16_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14680\,
            lcout => \spi_slave_1.miso_data_outZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_data_out_17_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14650\,
            lcout => \spi_slave_1.miso_data_outZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27495\,
            ce => \N__14551\,
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_out_10_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15189\,
            lcout => miso_data_in_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_11_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14973\,
            lcout => miso_data_in_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_12_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14769\,
            lcout => miso_data_in_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_13_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16590\,
            lcout => miso_data_in_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_14_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16386\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => miso_data_in_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_15_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16170\,
            lcout => miso_data_in_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_16_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18057\,
            lcout => miso_data_in_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.instr_out_17_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14674\,
            lcout => miso_data_in_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27499\,
            ce => \N__23994\,
            sr => \N__27124\
        );

    \sb_translator_1.addr_out_RNO_0_3_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14643\,
            in1 => \N__23009\,
            in2 => \_gnd_net_\,
            in3 => \N__14632\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_RNO_0_5_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23010\,
            in1 => \N__14604\,
            in2 => \_gnd_net_\,
            in3 => \N__14593\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIO2NL_0_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__19095\,
            in1 => \N__18966\,
            in2 => \N__19037\,
            in3 => \N__18994\,
            lcout => \sb_translator_1.state56_a_5_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16024\,
            lcout => \sb_translator_1.cnt19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27438\,
            ce => \N__22348\,
            sr => \N__27073\
        );

    \sb_translator_1.num_leds_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15997\,
            lcout => \sb_translator_1.num_ledsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27438\,
            ce => \N__22348\,
            sr => \N__27073\
        );

    \sb_translator_1.cnt_ram_read_RNIPFJ32_1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010101"
        )
    port map (
            in0 => \N__22405\,
            in1 => \N__17451\,
            in2 => \N__17418\,
            in3 => \N__22259\,
            lcout => \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_RNINT0G1_0_1_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__17447\,
            in1 => \N__17402\,
            in2 => \_gnd_net_\,
            in3 => \N__22401\,
            lcout => \sb_translator_1.send_leds_n_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_RNINT0G1_1_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__22403\,
            in1 => \_gnd_net_\,
            in2 => \N__17417\,
            in3 => \N__17450\,
            lcout => \sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_RNINT0G1_1_1_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17448\,
            in1 => \N__17406\,
            in2 => \_gnd_net_\,
            in3 => \N__22402\,
            lcout => \sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_RNINT0G1_2_1_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__22404\,
            in1 => \_gnd_net_\,
            in2 => \N__17416\,
            in3 => \N__17449\,
            lcout => \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIH2E91_9_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \N__20436\,
            in1 => \N__15923\,
            in2 => \N__15873\,
            in3 => \N__19181\,
            lcout => \sb_translator_1.num_leds_RNIH2E91Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIRUGT_10_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__15895\,
            in1 => \N__15868\,
            in2 => \_gnd_net_\,
            in3 => \N__19148\,
            lcout => \sb_translator_1.num_leds_RNIRUGTZ0Z_10\,
            ltout => \sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIP02R1_11_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20865\,
            in1 => \N__21387\,
            in2 => \N__14701\,
            in3 => \N__15894\,
            lcout => \sb_translator_1.num_leds_RNIP02R1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIU1HT_11_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__15896\,
            in1 => \_gnd_net_\,
            in2 => \N__21398\,
            in3 => \N__20866\,
            lcout => \sb_translator_1.num_leds_RNIU1HTZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIHKEQ_9_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__15867\,
            in1 => \N__15924\,
            in2 => \_gnd_net_\,
            in3 => \N__19180\,
            lcout => \sb_translator_1.num_leds_RNIHKEQZ0Z_9\,
            ltout => \sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNICJVN1_10_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__15893\,
            in1 => \N__15863\,
            in2 => \N__15844\,
            in3 => \N__19147\,
            lcout => \sb_translator_1.num_leds_RNICJVN1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI39BU_10_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19183\,
            lcout => \sb_translator_1.ram_sel_6_0_0_a2_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI39BU_0_10_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__19182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19149\,
            lcout => \sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__22203\,
            in2 => \_gnd_net_\,
            in3 => \N__18997\,
            lcout => addr_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22199\,
            in1 => \_gnd_net_\,
            in2 => \N__15571\,
            in3 => \N__18970\,
            lcout => addr_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_2_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18940\,
            in1 => \N__22204\,
            in2 => \_gnd_net_\,
            in3 => \N__15355\,
            lcout => addr_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22200\,
            in1 => \N__15139\,
            in2 => \_gnd_net_\,
            in3 => \N__18915\,
            lcout => addr_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_4_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22537\,
            in1 => \N__22205\,
            in2 => \_gnd_net_\,
            in3 => \N__18888\,
            lcout => addr_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_5_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22201\,
            in1 => \N__16759\,
            in2 => \_gnd_net_\,
            in3 => \N__18857\,
            lcout => addr_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_6_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22483\,
            in1 => \N__22206\,
            in2 => \_gnd_net_\,
            in3 => \N__18830\,
            lcout => addr_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.addr_out_7_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22202\,
            in1 => \_gnd_net_\,
            in2 => \N__22900\,
            in3 => \N__19244\,
            lcout => addr_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27452\,
            ce => \N__18027\,
            sr => \N__27080\
        );

    \sb_translator_1.cnt_RNILAHE_2_10_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17367\,
            in2 => \_gnd_net_\,
            in3 => \N__17319\,
            lcout => \sb_translator_1.cnt_RNILAHE_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI39BU_1_10_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__19185\,
            in1 => \N__19152\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI39BU_2_10_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19184\,
            in2 => \_gnd_net_\,
            in3 => \N__19153\,
            lcout => \sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_tmp_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16023\,
            in2 => \_gnd_net_\,
            in3 => \N__22015\,
            lcout => \sb_translator_1.instr_tmpZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27459\,
            ce => \N__16975\,
            sr => \N__27085\
        );

    \sb_translator_1.instr_tmp_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22013\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15996\,
            lcout => \sb_translator_1.instr_tmpZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27459\,
            ce => \N__16975\,
            sr => \N__27085\
        );

    \sb_translator_1.instr_tmp_2_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15957\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \sb_translator_1.instr_tmpZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27459\,
            ce => \N__16975\,
            sr => \N__27085\
        );

    \sb_translator_1.instr_tmp_3_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17025\,
            lcout => \sb_translator_1.instr_tmpZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27459\,
            ce => \N__16975\,
            sr => \N__27085\
        );

    \sb_translator_1.instr_tmp_4_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17001\,
            in2 => \_gnd_net_\,
            in3 => \N__22017\,
            lcout => \sb_translator_1.instr_tmpZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27459\,
            ce => \N__16975\,
            sr => \N__27085\
        );

    \sb_translator_1.rgb_data_tmp_18_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20994\,
            in1 => \N__21615\,
            in2 => \N__21576\,
            in3 => \N__21541\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27467\,
            ce => \N__25058\,
            sr => \N__27090\
        );

    \sb_translator_1.rgb_data_tmp_16_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20002\,
            in1 => \N__19940\,
            in2 => \N__19970\,
            in3 => \N__19895\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27467\,
            ce => \N__25058\,
            sr => \N__27090\
        );

    \sb_translator_1.ram_we_6_0_0_a2_1_7_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17629\,
            in1 => \N__17576\,
            in2 => \_gnd_net_\,
            in3 => \N__17681\,
            lcout => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_6_0_0_a2_2_11_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17682\,
            in1 => \N__17630\,
            in2 => \_gnd_net_\,
            in3 => \N__17577\,
            lcout => \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNIEL0N9_0_6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16888\,
            lcout => \sb_translator_1.state_RNIEL0N9_0Z0Z_6\,
            ltout => \sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNIOH7V9_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22009\,
            in2 => \N__16867\,
            in3 => \N__16863\,
            lcout => \sb_translator_1.state_RNIOH7V9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNI88IGA_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17493\,
            in2 => \_gnd_net_\,
            in3 => \N__17458\,
            lcout => \sb_translator_1.state_RNI88IGAZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000001"
        )
    port map (
            in0 => \N__27208\,
            in1 => \N__22421\,
            in2 => \N__17452\,
            in3 => \N__22306\,
            lcout => \sb_translator_1.cnt_ram_readZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27474\,
            ce => 'H',
            sr => \N__27096\
        );

    \sb_translator_1.cnt_ram_read_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__22422\,
            in1 => \N__17443\,
            in2 => \N__17419\,
            in3 => \N__17812\,
            lcout => \sb_translator_1.cnt_ram_readZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27474\,
            ce => 'H',
            sr => \N__27096\
        );

    \sb_translator_1.state_leds_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__27207\,
            in1 => \N__22305\,
            in2 => \N__17997\,
            in3 => \N__17833\,
            lcout => \sb_translator_1.state_ledsZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27474\,
            ce => 'H',
            sr => \N__27096\
        );

    \sb_translator_1.send_leds_n_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001100"
        )
    port map (
            in0 => \N__17832\,
            in1 => \N__22062\,
            in2 => \N__22210\,
            in3 => \N__27770\,
            lcout => send_leds_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27474\,
            ce => 'H',
            sr => \N__27096\
        );

    \ws2812.new_data_req_RNO_1_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__27769\,
            in1 => \N__25408\,
            in2 => \_gnd_net_\,
            in3 => \N__26905\,
            lcout => \ws2812.new_data_req_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_a3_4_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17380\,
            in2 => \_gnd_net_\,
            in3 => \N__23064\,
            lcout => \demux.N_422_i_0_a3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_RNILAHE_10_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17368\,
            in2 => \_gnd_net_\,
            in3 => \N__17320\,
            lcout => \sb_translator_1.ram_we_6_0_0_a2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_out_2_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20995\,
            in1 => \N__21604\,
            in2 => \N__21575\,
            in3 => \N__21539\,
            lcout => miso_data_in_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27483\,
            ce => \N__23992\,
            sr => \N__27102\
        );

    \sb_translator_1.state_RNI2IIJ_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17235\,
            in1 => \N__22785\,
            in2 => \_gnd_net_\,
            in3 => \N__17050\,
            lcout => \sb_translator_1.num_leds_1_sqmuxa\,
            ltout => \sb_translator_1.num_leds_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_ram_read_RNO_0_1_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27206\,
            in2 => \N__17836\,
            in3 => \N__17831\,
            lcout => \sb_translator_1.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.instr_out_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19971\,
            in1 => \N__19994\,
            in2 => \N__19908\,
            in3 => \N__19930\,
            lcout => miso_data_in_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27483\,
            ce => \N__23992\,
            sr => \N__27102\
        );

    \sb_translator_1.ram_sel_6_0_0_a2_2_5_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17590\,
            in1 => \N__17642\,
            in2 => \_gnd_net_\,
            in3 => \N__17695\,
            lcout => \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_sel_6_0_0_a2_3_13_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17693\,
            in1 => \N__17643\,
            in2 => \_gnd_net_\,
            in3 => \N__17588\,
            lcout => \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_6_0_0_a2_1_0_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17587\,
            in1 => \N__17641\,
            in2 => \_gnd_net_\,
            in3 => \N__17692\,
            lcout => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.ram_we_6_0_0_a2_1_3_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17694\,
            in1 => \N__17644\,
            in2 => \_gnd_net_\,
            in3 => \N__17589\,
            lcout => \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_13_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__18301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18322\,
            lcout => \demux.N_238\,
            ltout => \demux.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_17_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18273\,
            in2 => \N__17497\,
            in3 => \N__18246\,
            lcout => \demux.N_242\,
            ltout => \demux.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_34_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19840\,
            in2 => \N__17953\,
            in3 => \N__18356\,
            lcout => \demux.N_424_i_0_a2Z0Z_34\,
            ltout => \demux.N_424_i_0_a2Z0Z_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19810\,
            in1 => \N__20221\,
            in2 => \N__17950\,
            in3 => \N__19756\,
            lcout => \demux.N_424_i_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20319\,
            in1 => \N__20267\,
            in2 => \N__20365\,
            in3 => \N__19666\,
            lcout => \demux.N_424_i_0_aZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_11_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101001"
        )
    port map (
            in0 => \N__18357\,
            in1 => \N__18373\,
            in2 => \N__20227\,
            in3 => \N__17905\,
            lcout => \demux.N_424_i_0_o2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_3_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__18302\,
            in1 => \N__18286\,
            in2 => \N__18253\,
            in3 => \N__18323\,
            lcout => \demux.N_424_i_0_o2_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_11_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20222\,
            in1 => \N__19757\,
            in2 => \N__19818\,
            in3 => \N__19384\,
            lcout => \demux.N_424_i_0_a2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_1_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18251\,
            in1 => \N__19532\,
            in2 => \N__18285\,
            in3 => \N__18343\,
            lcout => \demux.N_424_i_0_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_38_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17904\,
            in1 => \N__19844\,
            in2 => \N__20226\,
            in3 => \N__18372\,
            lcout => \demux.N_916\,
            ltout => \demux.N_916_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_8_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__19569\,
            in1 => \N__17880\,
            in2 => \N__17860\,
            in3 => \N__17856\,
            lcout => \demux.N_424_i_0_a2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_10_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18303\,
            in1 => \N__18341\,
            in2 => \N__18328\,
            in3 => \N__19551\,
            lcout => \demux.N_424_i_0_a2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_9_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18252\,
            in1 => \N__19533\,
            in2 => \N__18284\,
            in3 => \N__18342\,
            lcout => \demux.N_424_i_0_a2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_37_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20217\,
            in1 => \N__18371\,
            in2 => \N__19848\,
            in3 => \N__18358\,
            lcout => \demux.N_915\,
            ltout => \demux.N_915_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_3_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19550\,
            in1 => \N__18324\,
            in2 => \N__18307\,
            in3 => \N__18304\,
            lcout => \demux.N_424_i_0_a2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_12_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18274\,
            in2 => \_gnd_net_\,
            in3 => \N__18250\,
            lcout => \demux.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_8_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21430\,
            in1 => \N__22198\,
            in2 => \_gnd_net_\,
            in3 => \N__19219\,
            lcout => addr_out_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27500\,
            ce => \N__18031\,
            sr => \N__27125\
        );

    \sb_translator_1.state_leds_RNIVONR_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22197\,
            in1 => \_gnd_net_\,
            in2 => \N__17998\,
            in3 => \N__22873\,
            lcout => \sb_translator_1.state_leds_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_leds_RNIGMAH_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17993\,
            in2 => \_gnd_net_\,
            in3 => \N__22196\,
            lcout => \sb_translator_1.state_leds_RNIGMAHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_13_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__17974\,
            in1 => \N__17968\,
            in2 => \_gnd_net_\,
            in3 => \N__18530\,
            lcout => \spi_slave_1.miso_RNOZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_6_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__18531\,
            in1 => \N__18616\,
            in2 => \_gnd_net_\,
            in3 => \N__18610\,
            lcout => \spi_slave_1.miso_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_14_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__18595\,
            in1 => \N__18589\,
            in2 => \_gnd_net_\,
            in3 => \N__18581\,
            lcout => OPEN,
            ltout => \spi_slave_1.N_58_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.miso_RNO_9_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__18532\,
            in1 => \_gnd_net_\,
            in2 => \N__18463\,
            in3 => \N__18460\,
            lcout => \spi_slave_1.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_1.mosi_data_out_15_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18442\,
            lcout => mosi_data_out_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27433\,
            ce => \N__18427\,
            sr => \N__27069\
        );

    \sb_translator_1.cnt_leds_RNI50UT_5_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101101001"
        )
    port map (
            in0 => \N__18405\,
            in1 => \N__18858\,
            in2 => \N__18655\,
            in3 => \N__20104\,
            lcout => \sb_translator_1.cnt_leds_RNI50UTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIK1VE_5_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18651\,
            in2 => \N__18862\,
            in3 => \N__18403\,
            lcout => \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5\,
            ltout => \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIB6UT_6_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18404\,
            in1 => \N__18832\,
            in2 => \N__18409\,
            in3 => \N__18800\,
            lcout => \sb_translator_1.cnt_leds_RNIB6UTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIN4VE_6_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010000"
        )
    port map (
            in0 => \N__18831\,
            in1 => \_gnd_net_\,
            in2 => \N__18804\,
            in3 => \N__18406\,
            lcout => \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6\,
            ltout => \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIHCUT_7_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18765\,
            in1 => \N__18796\,
            in2 => \N__18376\,
            in3 => \N__19245\,
            lcout => \sb_translator_1.cnt_leds_RNIHCUTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIQ7VE_7_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010000"
        )
    port map (
            in0 => \N__19246\,
            in1 => \_gnd_net_\,
            in2 => \N__18805\,
            in3 => \N__18763\,
            lcout => \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7\,
            ltout => \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNINIUT_8_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18764\,
            in1 => \N__18729\,
            in2 => \N__18769\,
            in3 => \N__19214\,
            lcout => \sb_translator_1.cnt_leds_RNINIUTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNITAVE_8_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011010100"
        )
    port map (
            in0 => \N__19215\,
            in1 => \N__18766\,
            in2 => \N__18733\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.cnt_leds_RNITAVEZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIO2NL_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101111010111"
        )
    port map (
            in0 => \N__19097\,
            in1 => \N__18968\,
            in2 => \N__19036\,
            in3 => \N__18995\,
            lcout => \sb_translator_1.N_318_i_i_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIBOUE_2_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__18938\,
            in1 => \N__19073\,
            in2 => \_gnd_net_\,
            in3 => \N__19023\,
            lcout => \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2\,
            ltout => \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIPJTT_3_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19075\,
            in1 => \N__18910\,
            in2 => \N__18691\,
            in3 => \N__18682\,
            lcout => \sb_translator_1.cnt_leds_RNIPJTTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIERUE_3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__18683\,
            in1 => \_gnd_net_\,
            in2 => \N__18916\,
            in3 => \N__19074\,
            lcout => \sb_translator_1.cnt_leds_RNIERUEZ0Z_3\,
            ltout => \sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIVPTT_4_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18650\,
            in1 => \N__18883\,
            in2 => \N__18688\,
            in3 => \N__18681\,
            lcout => \sb_translator_1.cnt_leds_RNIVPTTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIHUUE_4_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__18684\,
            in1 => \_gnd_net_\,
            in2 => \N__18889\,
            in3 => \N__18649\,
            lcout => \sb_translator_1.cnt_leds_RNIHUUEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI8LUE_1_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010110010"
        )
    port map (
            in0 => \N__19096\,
            in1 => \N__18967\,
            in2 => \N__19035\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.state56_a_5_44\,
            ltout => \sb_translator_1.state56_a_5_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIJDTT_2_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18937\,
            in1 => \N__19072\,
            in2 => \N__19045\,
            in3 => \N__19019\,
            lcout => \sb_translator_1.cnt_leds_RNIJDTTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22323\,
            in1 => \N__18996\,
            in2 => \_gnd_net_\,
            in3 => \N__18973\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \sb_translator_1.cnt_leds_cry_0\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22334\,
            in1 => \N__18969\,
            in2 => \_gnd_net_\,
            in3 => \N__18943\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_1\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_0\,
            carryout => \sb_translator_1.cnt_leds_cry_1\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22324\,
            in1 => \N__18939\,
            in2 => \_gnd_net_\,
            in3 => \N__18919\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_2\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_1\,
            carryout => \sb_translator_1.cnt_leds_cry_2\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_3_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22335\,
            in1 => \N__18914\,
            in2 => \_gnd_net_\,
            in3 => \N__18892\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_3\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_2\,
            carryout => \sb_translator_1.cnt_leds_cry_3\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_4_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22325\,
            in1 => \N__18887\,
            in2 => \_gnd_net_\,
            in3 => \N__18865\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_4\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_3\,
            carryout => \sb_translator_1.cnt_leds_cry_4\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_5_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22336\,
            in1 => \N__18856\,
            in2 => \_gnd_net_\,
            in3 => \N__18835\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_4\,
            carryout => \sb_translator_1.cnt_leds_cry_5\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_6_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22326\,
            in1 => \N__18829\,
            in2 => \_gnd_net_\,
            in3 => \N__18808\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_6\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_5\,
            carryout => \sb_translator_1.cnt_leds_cry_6\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_7_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22337\,
            in1 => \N__19243\,
            in2 => \_gnd_net_\,
            in3 => \N__19222\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_7\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_6\,
            carryout => \sb_translator_1.cnt_leds_cry_7\,
            clk => \N__27453\,
            ce => \N__19355\,
            sr => \N__27081\
        );

    \sb_translator_1.cnt_leds_8_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22333\,
            in1 => \N__19213\,
            in2 => \_gnd_net_\,
            in3 => \N__19192\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \sb_translator_1.cnt_leds_cry_8\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_9_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22321\,
            in1 => \N__21352\,
            in2 => \_gnd_net_\,
            in3 => \N__19189\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_9\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_8\,
            carryout => \sb_translator_1.cnt_leds_cry_9\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_10_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__19186\,
            in2 => \_gnd_net_\,
            in3 => \N__19156\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_10\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_9\,
            carryout => \sb_translator_1.cnt_leds_cry_10\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_11_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22318\,
            in1 => \N__19151\,
            in2 => \_gnd_net_\,
            in3 => \N__19120\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_11\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_10\,
            carryout => \sb_translator_1.cnt_leds_cry_11\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_12_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22331\,
            in1 => \N__21391\,
            in2 => \_gnd_net_\,
            in3 => \N__19117\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_12\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_11\,
            carryout => \sb_translator_1.cnt_leds_cry_12\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_13_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22319\,
            in1 => \N__20842\,
            in2 => \_gnd_net_\,
            in3 => \N__19114\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_13\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_12\,
            carryout => \sb_translator_1.cnt_leds_cry_13\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_14_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22332\,
            in1 => \N__20743\,
            in2 => \_gnd_net_\,
            in3 => \N__19111\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_14\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_13\,
            carryout => \sb_translator_1.cnt_leds_cry_14\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_15_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22320\,
            in1 => \N__20905\,
            in2 => \_gnd_net_\,
            in3 => \N__19372\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_15\,
            ltout => OPEN,
            carryin => \sb_translator_1.cnt_leds_cry_14\,
            carryout => \sb_translator_1.cnt_leds_cry_15\,
            clk => \N__27460\,
            ce => \N__19366\,
            sr => \N__27086\
        );

    \sb_translator_1.cnt_leds_16_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__20599\,
            in1 => \N__22322\,
            in2 => \_gnd_net_\,
            in3 => \N__19369\,
            lcout => \sb_translator_1.cnt_ledsZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27468\,
            ce => \N__19365\,
            sr => \N__27091\
        );

    \sb_translator_1.rgb_data_tmp_2_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20980\,
            in1 => \N__21619\,
            in2 => \N__21574\,
            in3 => \N__21538\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27475\,
            ce => \N__25430\,
            sr => \N__27097\
        );

    \demux.N_424_i_0_a3_4_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__23073\,
            lcout => \demux.N_424_i_0_a3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__19327\,
            in1 => \N__23371\,
            in2 => \_gnd_net_\,
            in3 => \N__20644\,
            lcout => OPEN,
            ltout => \demux.N_424_i_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_7_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__19309\,
            in2 => \N__19294\,
            in3 => \N__23302\,
            lcout => \demux.N_424_i_0_o2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19291\,
            in2 => \_gnd_net_\,
            in3 => \N__25836\,
            lcout => \demux.N_424_i_0_aZ0Z3\,
            ltout => \demux.N_424_i_0_aZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20001\,
            in1 => \N__19947\,
            in2 => \N__19276\,
            in3 => \N__19894\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27475\,
            ce => \N__25430\,
            sr => \N__27097\
        );

    \demux.N_421_i_0_o2_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23477\,
            in1 => \N__19273\,
            in2 => \N__19261\,
            in3 => \N__23408\,
            lcout => OPEN,
            ltout => \demux.N_421_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__19519\,
            in1 => \N__23367\,
            in2 => \N__19507\,
            in3 => \N__19390\,
            lcout => \demux.N_421_i_0_o2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_a3_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19504\,
            lcout => \demux.N_422_i_0_aZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__19489\,
            in1 => \N__19477\,
            in2 => \N__23424\,
            in3 => \N__23478\,
            lcout => OPEN,
            ltout => \demux.N_422_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__23368\,
            in1 => \_gnd_net_\,
            in2 => \N__19465\,
            in3 => \N__19462\,
            lcout => OPEN,
            ltout => \demux.N_422_i_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_7_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19450\,
            in1 => \N__19444\,
            in2 => \N__19432\,
            in3 => \N__23298\,
            lcout => \demux.N_422_i_0_o2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_a3_5_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23297\,
            in2 => \_gnd_net_\,
            in3 => \N__19429\,
            lcout => OPEN,
            ltout => \demux.N_423_i_0_a3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__19417\,
            in1 => \N__23346\,
            in2 => \N__19405\,
            in3 => \N__19672\,
            lcout => \demux.N_423_i_0_o2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_a3_4_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23055\,
            in2 => \_gnd_net_\,
            in3 => \N__19402\,
            lcout => \demux.N_837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_12_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__19817\,
            in1 => \N__19767\,
            in2 => \_gnd_net_\,
            in3 => \N__19383\,
            lcout => \demux.N_918\,
            ltout => \demux.N_918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_5_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20316\,
            in1 => \N__20361\,
            in2 => \N__19705\,
            in3 => \N__20274\,
            lcout => \demux.N_424_i_0_a2Z0Z_5\,
            ltout => \demux.N_424_i_0_a2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_0_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__23452\,
            in1 => \N__19702\,
            in2 => \N__19690\,
            in3 => \N__19687\,
            lcout => \demux.N_423_i_0_o2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_7_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20318\,
            in1 => \N__20359\,
            in2 => \N__20275\,
            in3 => \N__19665\,
            lcout => \demux.N_424_i_0_a2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_44_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20360\,
            in1 => \N__20273\,
            in2 => \_gnd_net_\,
            in3 => \N__20317\,
            lcout => \demux.N_917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_13_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25848\,
            in1 => \N__25747\,
            in2 => \N__25723\,
            in3 => \N__25655\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27496\,
            ce => \N__21503\,
            sr => \N__27115\
        );

    \sb_translator_1.rgb_data_tmp_11_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24220\,
            in1 => \N__25849\,
            in2 => \N__24263\,
            in3 => \N__24177\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27496\,
            ce => \N__21503\,
            sr => \N__27115\
        );

    \demux.N_424_i_0_o2_0_8_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__19615\,
            in1 => \N__19603\,
            in2 => \_gnd_net_\,
            in3 => \N__19576\,
            lcout => OPEN,
            ltout => \demux.N_424_i_0_o2_0_8Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_8_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__19558\,
            in1 => \N__19552\,
            in2 => \N__19537\,
            in3 => \N__19534\,
            lcout => OPEN,
            ltout => \demux.N_424_i_0_o2_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19729\,
            in1 => \N__20062\,
            in2 => \N__20056\,
            in3 => \N__20053\,
            lcout => \demux.N_424_i_0_o2Z0Z_0\,
            ltout => \demux.N_424_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__24092\,
            in1 => \N__24121\,
            in2 => \N__20047\,
            in3 => \N__24044\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27496\,
            ce => \N__21503\,
            sr => \N__27115\
        );

    \demux.N_424_i_0_o2_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__20044\,
            in1 => \N__24478\,
            in2 => \N__20032\,
            in3 => \N__24411\,
            lcout => OPEN,
            ltout => \demux.N_424_i_0_o2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_8_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24326\,
            in1 => \N__20017\,
            in2 => \N__20005\,
            in3 => \N__19858\,
            lcout => \demux.N_424_i_0_o2Z0Z_8\,
            ltout => \demux.N_424_i_0_o2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_8_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19975\,
            in1 => \N__19948\,
            in2 => \N__19912\,
            in3 => \N__19909\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27501\,
            ce => \N__21517\,
            sr => \N__27126\
        );

    \demux.N_424_i_0_a3_7_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19876\,
            lcout => \demux.N_424_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_a2_33_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20269\,
            in1 => \_gnd_net_\,
            in2 => \N__20320\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \demux.N_906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__19819\,
            in2 => \N__19771\,
            in3 => \N__19768\,
            lcout => \demux.N_424_i_0_o2_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_a3_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19723\,
            in2 => \_gnd_net_\,
            in3 => \N__23930\,
            lcout => \demux.N_420_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_15_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20358\,
            in1 => \N__20312\,
            in2 => \_gnd_net_\,
            in3 => \N__20268\,
            lcout => \demux.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_a3_7_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23922\,
            in2 => \_gnd_net_\,
            in3 => \N__20197\,
            lcout => \demux.N_419_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_0_c_THRU_CRY_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20172\,
            in2 => \N__20179\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \sb_translator_1.state56_a_5_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIJ5J22_0_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20158\,
            in2 => \N__20152\,
            in3 => \N__20143\,
            lcout => \sb_translator_1.state56_a_5_2\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_0_c_THRU_CO\,
            carryout => \sb_translator_1.state56_a_5_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_0_c_RNIUH4N1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20140\,
            in2 => \N__20134\,
            in3 => \N__20125\,
            lcout => \sb_translator_1.state56_a_5_3\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_0\,
            carryout => \sb_translator_1.state56_a_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_1_c_RNI8T5N1_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20122\,
            in2 => \N__20116\,
            in3 => \N__20107\,
            lcout => \sb_translator_1.state56_a_5_4\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_1\,
            carryout => \sb_translator_1.state56_a_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_2_c_RNII87N1_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20103\,
            in2 => \N__20092\,
            in3 => \N__20083\,
            lcout => \sb_translator_1.state56_a_5_5\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_2\,
            carryout => \sb_translator_1.state56_a_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_3_c_RNISJ8N1_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20080\,
            in2 => \N__20074\,
            in3 => \N__20065\,
            lcout => \sb_translator_1.state56_a_5_6\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_3\,
            carryout => \sb_translator_1.state56_a_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_4_c_RNI6V9N1_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20521\,
            in2 => \N__20515\,
            in3 => \N__20506\,
            lcout => \sb_translator_1.state56_a_5_7\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_4\,
            carryout => \sb_translator_1.state56_a_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_5_c_RNIGABN1_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20503\,
            in2 => \N__20497\,
            in3 => \N__20488\,
            lcout => \sb_translator_1.state56_a_5_8\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_5\,
            carryout => \sb_translator_1.state56_a_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_6_c_RNIQLCN1_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20485\,
            in2 => \N__20475\,
            in3 => \N__20452\,
            lcout => \sb_translator_1.state56_a_5_9\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \sb_translator_1.state56_a_5_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_7_c_RNII4T22_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \N__20440\,
            in3 => \N__20422\,
            lcout => \sb_translator_1.state56_a_5_10\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_7\,
            carryout => \sb_translator_1.state56_a_5_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_8_c_RNIVTUS2_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20419\,
            in2 => \N__20410\,
            in3 => \N__20398\,
            lcout => \sb_translator_1.state56_a_5_11\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_8\,
            carryout => \sb_translator_1.state56_a_5_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_9_c_RNINN433_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20395\,
            in2 => \N__20386\,
            in3 => \N__20374\,
            lcout => \sb_translator_1.state56_a_5_12\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_9\,
            carryout => \sb_translator_1.state56_a_5_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_10_c_RNI8BIQ2_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20554\,
            in2 => \N__20574\,
            in3 => \N__20371\,
            lcout => \sb_translator_1.state56_a_5_13\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_10\,
            carryout => \sb_translator_1.state56_a_5_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_11_c_RNIIMJQ2_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20827\,
            in2 => \N__20728\,
            in3 => \N__20368\,
            lcout => \sb_translator_1.state56_a_5_14\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_11\,
            carryout => \sb_translator_1.state56_a_5_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_12_c_RNIS1LQ2_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20530\,
            in2 => \N__20545\,
            in3 => \N__20608\,
            lcout => \sb_translator_1.state56_a_5_15\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_12\,
            carryout => \sb_translator_1.state56_a_5_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_13_c_RNIK1552_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20584\,
            in2 => \N__20890\,
            in3 => \N__20605\,
            lcout => \sb_translator_1.state56_a_5_16\,
            ltout => OPEN,
            carryin => \sb_translator_1.state56_a_5_cry_13\,
            carryout => \sb_translator_1.state56_a_5_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_14_c_RNI7UEO_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20916\,
            in1 => \N__20949\,
            in2 => \_gnd_net_\,
            in3 => \N__20602\,
            lcout => \sb_translator_1.state56_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_15_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22945\,
            lcout => \sb_translator_1.num_ledsZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27469\,
            ce => \N__22355\,
            sr => \N__27092\
        );

    \sb_translator_1.cnt_leds_RNI7Q5F_16_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20598\,
            lcout => \sb_translator_1.cnt_leds_i_16\,
            ltout => \sb_translator_1.cnt_leds_i_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.num_leds_RNIOJBM_15_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__20947\,
            in1 => \_gnd_net_\,
            in2 => \N__20587\,
            in3 => \_gnd_net_\,
            lcout => \sb_translator_1.num_leds_RNIOJBMZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIV62R1_13_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \N__20575\,
            in1 => \N__20877\,
            in2 => \N__20782\,
            in3 => \N__20840\,
            lcout => \sb_translator_1.cnt_leds_RNIV62R1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI48HT_14_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__20812\,
            in1 => \N__20781\,
            in2 => \_gnd_net_\,
            in3 => \N__20742\,
            lcout => \sb_translator_1.cnt_leds_RNI48HTZ0Z_14\,
            ltout => \sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIBJ2R1_15_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20903\,
            in1 => \N__20946\,
            in2 => \N__20533\,
            in3 => \N__20814\,
            lcout => \sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNIE5NC1_15_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__20815\,
            in1 => \N__20948\,
            in2 => \N__20920\,
            in3 => \N__20904\,
            lcout => \sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI15HT_13_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__20780\,
            in1 => \N__20878\,
            in2 => \_gnd_net_\,
            in3 => \N__20841\,
            lcout => \sb_translator_1.cnt_leds_RNI15HTZ0Z_13\,
            ltout => \sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI5D2R1_14_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20813\,
            in1 => \N__20776\,
            in2 => \N__20746\,
            in3 => \N__20741\,
            lcout => \sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_8_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__23809\,
            in1 => \N__24361\,
            in2 => \N__20716\,
            in3 => \N__21268\,
            lcout => \demux.N_422_i_0_o2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20701\,
            in1 => \N__24435\,
            in2 => \N__20686\,
            in3 => \N__23956\,
            lcout => \demux.N_418_i_0_o2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_424_i_0_o2_0_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23479\,
            in1 => \N__20674\,
            in2 => \N__20659\,
            in3 => \N__23412\,
            lcout => \demux.N_424_i_0_o2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_a3_4_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20638\,
            in2 => \_gnd_net_\,
            in3 => \N__23074\,
            lcout => \demux.N_420_i_0_a3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_a3_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20623\,
            in2 => \_gnd_net_\,
            in3 => \N__24505\,
            lcout => OPEN,
            ltout => \demux.N_884_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_8_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__21154\,
            in1 => \N__21148\,
            in2 => \N__21133\,
            in3 => \N__21073\,
            lcout => \demux.N_418_i_0_o2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_a3_7_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23951\,
            in2 => \_gnd_net_\,
            in3 => \N__21130\,
            lcout => \demux.N_421_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21115\,
            in1 => \N__24504\,
            in2 => \N__21100\,
            in3 => \N__24434\,
            lcout => OPEN,
            ltout => \demux.N_421_i_0_o2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_8_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21088\,
            in1 => \N__21072\,
            in2 => \N__21025\,
            in3 => \N__21022\,
            lcout => OPEN,
            ltout => \demux.N_421_i_0_o2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_421_i_0_o2_10_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21016\,
            in1 => \N__23296\,
            in2 => \N__21004\,
            in3 => \N__21001\,
            lcout => \demux.N_421_i_0_o2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_15_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23714\,
            in1 => \N__23884\,
            in2 => \N__23700\,
            in3 => \N__23771\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27497\,
            ce => \N__21516\,
            sr => \N__27116\
        );

    \sb_translator_1.rgb_data_tmp_14_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23617\,
            in1 => \N__23645\,
            in2 => \N__23588\,
            in3 => \N__23558\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27497\,
            ce => \N__21516\,
            sr => \N__27116\
        );

    \sb_translator_1.rgb_data_tmp_12_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25623\,
            in1 => \N__25574\,
            in2 => \N__25539\,
            in3 => \N__25477\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27497\,
            ce => \N__21516\,
            sr => \N__27116\
        );

    \sb_translator_1.rgb_data_tmp_10_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20990\,
            in1 => \N__21614\,
            in2 => \N__21583\,
            in3 => \N__21540\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27497\,
            ce => \N__21516\,
            sr => \N__27116\
        );

    \sb_translator_1.addr_out_RNO_0_8_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23008\,
            in1 => \N__21469\,
            in2 => \_gnd_net_\,
            in3 => \N__21457\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.cnt_leds_RNI1VFQ_2_9_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21997\,
            in1 => \N__21416\,
            in2 => \_gnd_net_\,
            in3 => \N__21363\,
            lcout => \sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_a3_7_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__23950\,
            in1 => \_gnd_net_\,
            in2 => \N__21283\,
            in3 => \_gnd_net_\,
            lcout => \demux.N_422_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_7_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23295\,
            in1 => \N__21259\,
            in2 => \N__21739\,
            in3 => \N__21760\,
            lcout => \demux.N_417_i_0_o2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_a3_7_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23949\,
            in2 => \_gnd_net_\,
            in3 => \N__21247\,
            lcout => \demux.N_423_i_0_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21229\,
            in1 => \N__24506\,
            in2 => \N__21217\,
            in3 => \N__24436\,
            lcout => OPEN,
            ltout => \demux.N_423_i_0_o2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_8_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21202\,
            in1 => \N__24354\,
            in2 => \N__21187\,
            in3 => \N__21184\,
            lcout => OPEN,
            ltout => \demux.N_423_i_0_o2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_423_i_0_o2_10_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21178\,
            in1 => \N__23072\,
            in2 => \N__21163\,
            in3 => \N__21160\,
            lcout => \demux.N_423_i_0_o2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__23480\,
            in1 => \N__21808\,
            in2 => \N__23425\,
            in3 => \N__21796\,
            lcout => OPEN,
            ltout => \demux.N_417_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21778\,
            in2 => \N__21763\,
            in3 => \N__23369\,
            lcout => \demux.N_417_i_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_a3_4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21754\,
            in2 => \_gnd_net_\,
            in3 => \N__23056\,
            lcout => \demux.N_417_i_0_a3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__23481\,
            in1 => \N__21730\,
            in2 => \N__23426\,
            in3 => \N__21718\,
            lcout => OPEN,
            ltout => \demux.N_419_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21700\,
            in1 => \N__23370\,
            in2 => \N__21685\,
            in3 => \N__21655\,
            lcout => OPEN,
            ltout => \demux.N_419_i_0_o2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_10_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23057\,
            in1 => \N__21682\,
            in2 => \N__21667\,
            in3 => \N__21625\,
            lcout => \demux.N_419_i_0_o2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_a3_5_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23272\,
            in2 => \_gnd_net_\,
            in3 => \N__21664\,
            lcout => \demux.N_419_i_0_a3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_8_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__24353\,
            in1 => \N__24526\,
            in2 => \N__21649\,
            in3 => \N__21631\,
            lcout => \demux.N_419_i_0_o2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_2_c_RNILP7UD_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__22471\,
            in1 => \N__22465\,
            in2 => \N__22459\,
            in3 => \N__22105\,
            lcout => OPEN,
            ltout => \sb_translator_1.N_318_i_i_o2_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_10_c_RNIMPSBK_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__22450\,
            in1 => \N__22444\,
            in2 => \N__22438\,
            in3 => \N__22435\,
            lcout => OPEN,
            ltout => \sb_translator_1.N_318_i_i_o2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_RNI41J131_7_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110110011"
        )
    port map (
            in0 => \N__22151\,
            in1 => \N__22426\,
            in2 => \N__22369\,
            in3 => \N__22834\,
            lcout => \sb_translator_1.N_712\,
            ltout => \sb_translator_1.N_712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_7_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22366\,
            in3 => \N__22347\,
            lcout => \sb_translator_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27461\,
            ce => 'H',
            sr => \N__27087\
        );

    \sb_translator_1.cnt_leds_RNI8VOI7_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22135\,
            in1 => \N__22129\,
            in2 => \N__22123\,
            in3 => \N__22111\,
            lcout => \sb_translator_1.N_318_i_i_o2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22099\,
            in1 => \N__21856\,
            in2 => \N__22828\,
            in3 => \N__22081\,
            lcout => \sb_translator_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27461\,
            ce => 'H',
            sr => \N__27087\
        );

    \sb_translator_1.state_6_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__22821\,
            in1 => \N__22752\,
            in2 => \N__22645\,
            in3 => \N__21855\,
            lcout => \sb_translator_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27470\,
            ce => 'H',
            sr => \N__27093\
        );

    \sb_translator_1.state56_a_5_cry_13_c_RNICLCM7_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21835\,
            in1 => \N__21829\,
            in2 => \N__21823\,
            in3 => \N__21814\,
            lcout => OPEN,
            ltout => \sb_translator_1.N_318_i_i_o2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state56_a_5_cry_12_c_RNIINPVD_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22855\,
            in1 => \N__22849\,
            in2 => \N__22843\,
            in3 => \N__22840\,
            lcout => \sb_translator_1.N_318_i_i_o2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.state_1_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__22639\,
            in1 => \_gnd_net_\,
            in2 => \N__22784\,
            in3 => \N__22820\,
            lcout => \sb_translator_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27470\,
            ce => 'H',
            sr => \N__27093\
        );

    \sb_translator_1.state_ns_i_i_0_0_o3_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22751\,
            in2 => \_gnd_net_\,
            in3 => \N__22638\,
            lcout => \sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_3_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__27750\,
            in1 => \N__27864\,
            in2 => \N__27607\,
            in3 => \N__26473\,
            lcout => \ws2812.rgb_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27476\,
            ce => 'H',
            sr => \N__27098\
        );

    \ws2812.rgb_counter_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000010001"
        )
    port map (
            in0 => \N__27862\,
            in1 => \N__27749\,
            in2 => \_gnd_net_\,
            in3 => \N__27911\,
            lcout => \ws2812.rgb_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27476\,
            ce => 'H',
            sr => \N__27098\
        );

    \ws2812.bit_counter_0_1_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__27574\,
            in1 => \N__27863\,
            in2 => \_gnd_net_\,
            in3 => \N__24721\,
            lcout => \ws2812.bit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27476\,
            ce => 'H',
            sr => \N__27098\
        );

    \sb_translator_1.addr_out_RNO_0_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22582\,
            in1 => \N__22978\,
            in2 => \_gnd_net_\,
            in3 => \N__22564\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_RNO_0_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22525\,
            in1 => \N__22507\,
            in2 => \_gnd_net_\,
            in3 => \N__22979\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.addr_out_RNO_0_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22980\,
            in1 => \N__22944\,
            in2 => \_gnd_net_\,
            in3 => \N__22926\,
            lcout => \sb_translator_1.addr_out_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNING643_4_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__25400\,
            in1 => \N__26407\,
            in2 => \N__27747\,
            in3 => \N__26898\,
            lcout => \ws2812.bit_counter_0_RNING643Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNO_0_5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100001011010"
        )
    port map (
            in0 => \N__26899\,
            in1 => \N__27723\,
            in2 => \N__25231\,
            in3 => \N__25401\,
            lcout => \ws2812.un1_bit_counter_12_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNI6OQB3_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__25396\,
            in1 => \N__24664\,
            in2 => \N__27745\,
            in3 => \N__26894\,
            lcout => \ws2812.bit_counter_RNI6OQB3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNI7PQB3_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__26895\,
            in1 => \N__27715\,
            in2 => \N__24619\,
            in3 => \N__25397\,
            lcout => \ws2812.bit_counter_RNI7PQB3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNI8QQB3_4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__25399\,
            in1 => \N__24838\,
            in2 => \N__27746\,
            in3 => \N__26896\,
            lcout => \ws2812.bit_counter_RNI8QQB3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNI9RQB3_5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__26897\,
            in1 => \N__27719\,
            in2 => \N__26368\,
            in3 => \N__25398\,
            lcout => \ws2812.bit_counter_RNI9RQB3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.new_data_req_RNO_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__25402\,
            in1 => \N__27600\,
            in2 => \N__27748\,
            in3 => \N__26900\,
            lcout => OPEN,
            ltout => \ws2812.N_140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.new_data_req_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101100"
        )
    port map (
            in0 => \N__22888\,
            in1 => \N__22869\,
            in2 => \N__22876\,
            in3 => \N__25403\,
            lcout => ws2812_next_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27484\,
            ce => 'H',
            sr => \N__27103\
        );

    \sb_translator_1.rgb_data_out_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23182\,
            lcout => rgb_data_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \sb_translator_1.rgb_data_out_10_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_data_out_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \sb_translator_1.rgb_data_out_12_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23164\,
            lcout => rgb_data_out_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \sb_translator_1.rgb_data_out_18_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23155\,
            lcout => rgb_data_out_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \sb_translator_1.rgb_data_out_15_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23146\,
            lcout => rgb_data_out_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \sb_translator_1.rgb_data_out_16_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => rgb_data_out_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27490\,
            ce => \N__27193\,
            sr => \N__27111\
        );

    \demux.N_418_i_0_o2_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23125\,
            in1 => \N__23365\,
            in2 => \N__23434\,
            in3 => \N__23116\,
            lcout => OPEN,
            ltout => \demux.N_418_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__23488\,
            in1 => \_gnd_net_\,
            in2 => \N__23110\,
            in3 => \N__23107\,
            lcout => OPEN,
            ltout => \demux.N_418_i_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_o2_7_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__23089\,
            in1 => \N__23512\,
            in2 => \N__23077\,
            in3 => \N__23071\,
            lcout => \demux.N_418_i_0_o2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_418_i_0_a3_5_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23524\,
            in2 => \_gnd_net_\,
            in3 => \N__23293\,
            lcout => \demux.N_880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23506\,
            in1 => \N__23487\,
            in2 => \N__23433\,
            in3 => \N__23377\,
            lcout => OPEN,
            ltout => \demux.N_420_i_0_o2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__23366\,
            in1 => \_gnd_net_\,
            in2 => \N__23317\,
            in3 => \N__23314\,
            lcout => OPEN,
            ltout => \demux.N_420_i_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23294\,
            in1 => \N__23236\,
            in2 => \N__23221\,
            in3 => \N__23218\,
            lcout => \demux.N_420_i_0_o2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_a3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23209\,
            in2 => \_gnd_net_\,
            in3 => \N__25854\,
            lcout => \demux.N_888\,
            ltout => \demux.N_888_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_7_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23883\,
            in1 => \N__23779\,
            in2 => \N__23197\,
            in3 => \N__23699\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27502\,
            ce => \N__25437\,
            sr => \N__27127\
        );

    \sb_translator_1.rgb_data_tmp_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25859\,
            in1 => \N__24256\,
            in2 => \N__24218\,
            in3 => \N__24172\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27502\,
            ce => \N__25437\,
            sr => \N__27127\
        );

    \sb_translator_1.rgb_data_tmp_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25855\,
            in1 => \N__24131\,
            in2 => \N__24085\,
            in3 => \N__24046\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27502\,
            ce => \N__25437\,
            sr => \N__27127\
        );

    \demux.N_418_i_0_a3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23194\,
            in2 => \_gnd_net_\,
            in3 => \N__25852\,
            lcout => \demux.N_874\,
            ltout => \demux.N_874_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__23582\,
            in2 => \N__23797\,
            in3 => \N__23551\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27502\,
            ce => \N__25437\,
            sr => \N__27127\
        );

    \demux.N_420_i_0_a3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23794\,
            in2 => \_gnd_net_\,
            in3 => \N__25853\,
            lcout => \demux.N_420_i_0_aZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_tmp_23_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23721\,
            in1 => \N__23882\,
            in2 => \N__23701\,
            in3 => \N__23770\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27507\,
            ce => \N__25077\,
            sr => \N__27130\
        );

    \sb_translator_1.rgb_data_tmp_22_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23625\,
            in1 => \N__23595\,
            in2 => \N__23658\,
            in3 => \N__23559\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27507\,
            ce => \N__25077\,
            sr => \N__27130\
        );

    \sb_translator_1.rgb_data_tmp_21_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25850\,
            in1 => \N__25757\,
            in2 => \N__25715\,
            in3 => \N__25656\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27507\,
            ce => \N__25077\,
            sr => \N__27130\
        );

    \sb_translator_1.rgb_data_tmp_19_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__24264\,
            in2 => \N__25867\,
            in3 => \N__24176\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27507\,
            ce => \N__25077\,
            sr => \N__27130\
        );

    \sb_translator_1.rgb_data_tmp_17_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24093\,
            in1 => \N__25851\,
            in2 => \N__24136\,
            in3 => \N__24043\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27507\,
            ce => \N__25077\,
            sr => \N__27130\
        );

    \sb_translator_1.instr_out_7_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23881\,
            in1 => \N__23778\,
            in2 => \N__23725\,
            in3 => \N__23698\,
            lcout => miso_data_in_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \sb_translator_1.instr_out_6_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23659\,
            in1 => \N__23629\,
            in2 => \N__23599\,
            in3 => \N__23560\,
            lcout => miso_data_in_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \sb_translator_1.instr_out_5_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25861\,
            in1 => \N__25765\,
            in2 => \N__25711\,
            in3 => \N__25654\,
            lcout => miso_data_in_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \sb_translator_1.instr_out_3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__24265\,
            in1 => \N__24219\,
            in2 => \N__24178\,
            in3 => \N__25862\,
            lcout => miso_data_in_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \sb_translator_1.instr_out_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25860\,
            in1 => \N__24135\,
            in2 => \N__24097\,
            in3 => \N__24045\,
            lcout => miso_data_in_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \sb_translator_1.instr_out_4_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25603\,
            in1 => \N__25581\,
            in2 => \N__25540\,
            in3 => \N__25484\,
            lcout => miso_data_in_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27511\,
            ce => \N__23991\,
            sr => \N__27134\
        );

    \demux.N_417_i_0_a3_7_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23971\,
            in2 => \_gnd_net_\,
            in3 => \N__23955\,
            lcout => OPEN,
            ltout => \demux.N_417_i_0_a3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_8_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__23899\,
            in1 => \N__23839\,
            in2 => \N__23887\,
            in3 => \N__24358\,
            lcout => \demux.N_417_i_0_o2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_417_i_0_o2_4_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24432\,
            in1 => \N__23857\,
            in2 => \N__24508\,
            in3 => \N__23845\,
            lcout => \demux.N_417_i_0_o2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_422_i_0_o2_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23833\,
            in1 => \N__24502\,
            in2 => \N__23824\,
            in3 => \N__24431\,
            lcout => \demux.N_422_i_0_o2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_419_i_0_o2_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__24430\,
            in1 => \N__24544\,
            in2 => \N__24507\,
            in3 => \N__24532\,
            lcout => \demux.N_419_i_0_o2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24520\,
            in1 => \N__24503\,
            in2 => \N__24451\,
            in3 => \N__24433\,
            lcout => OPEN,
            ltout => \demux.N_420_i_0_o2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \demux.N_420_i_0_o2_8_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24376\,
            in1 => \N__24359\,
            in2 => \N__24292\,
            in3 => \N__24289\,
            lcout => \demux.N_420_i_0_o2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIKD643_1_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__27734\,
            in1 => \N__26860\,
            in2 => \N__24769\,
            in3 => \N__25360\,
            lcout => \ws2812.bit_counter_0_RNIKD643Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNILE643_2_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001010"
        )
    port map (
            in0 => \N__26861\,
            in1 => \N__24895\,
            in2 => \N__25393\,
            in3 => \N__27735\,
            lcout => \ws2812.bit_counter_0_RNILE643Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIMF643_3_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__27736\,
            in1 => \N__25361\,
            in2 => \N__24868\,
            in3 => \N__26862\,
            lcout => \ws2812.bit_counter_0_RNIMF643Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.state_1_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__26863\,
            in1 => \N__27786\,
            in2 => \N__25394\,
            in3 => \N__27737\,
            lcout => \ws2812.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27471\,
            ce => 'H',
            sr => \N__27094\
        );

    \ws2812.un1_bit_counter_12_cry_0_c_RNO_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__27732\,
            in1 => \N__25355\,
            in2 => \N__25275\,
            in3 => \N__26858\,
            lcout => \ws2812.un1_bit_counter_12_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNI5NQB3_1_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__27733\,
            in1 => \N__26859\,
            in2 => \N__25303\,
            in3 => \N__25356\,
            lcout => \ws2812.bit_counter_RNI5NQB3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNIENHA_3_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24607\,
            lcout => \ws2812.un6_data_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIQAT2_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25181\,
            lcout => \ws2812.bit_counter_0_RNIQAT2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIRBT2_1_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24765\,
            lcout => \ws2812.bit_counter_0_RNIRBT2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIG4UQ_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24764\,
            in1 => \N__24655\,
            in2 => \N__24612\,
            in3 => \N__25180\,
            lcout => \ws2812.state_ns_0_i_o2_6_0\,
            ltout => \ws2812.state_ns_0_i_o2_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNISPQG2_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25311\,
            in2 => \N__24568\,
            in3 => \N__24906\,
            lcout => \ws2812.N_105\,
            ltout => \ws2812.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIJC643_0_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010110000"
        )
    port map (
            in0 => \N__27741\,
            in1 => \N__25369\,
            in2 => \N__24565\,
            in3 => \N__25182\,
            lcout => \ws2812.bit_counter_0_RNIJC643Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.state_RNIBU1P2_1_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24562\,
            in1 => \N__25312\,
            in2 => \N__25395\,
            in3 => \N__24907\,
            lcout => \ws2812.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNIDMHA_2_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24656\,
            lcout => \ws2812.un6_data_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un1_bit_counter_12_cry_0_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25270\,
            in2 => \N__24556\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \ws2812.un1_bit_counter_12_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25296\,
            in2 => \N__24793\,
            in3 => \N__24781\,
            lcout => \ws2812.bit_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_0\,
            carryout => \ws2812.un1_bit_counter_12_cry_1\,
            clk => \N__27485\,
            ce => 'H',
            sr => \N__27108\
        );

    \ws2812.bit_counter_0_RNO_0_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24778\,
            in2 => \N__25189\,
            in3 => \N__24772\,
            lcout => \ws2812.bit_counter_0_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_1\,
            carryout => \ws2812.un1_bit_counter_12_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNO_0_1_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24760\,
            in2 => \N__24733\,
            in3 => \N__24712\,
            lcout => \ws2812.bit_counter_0_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_2\,
            carryout => \ws2812.un1_bit_counter_12_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_2_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__27828\,
            in1 => \N__24889\,
            in2 => \N__24709\,
            in3 => \N__24697\,
            lcout => \ws2812.bit_counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_3\,
            carryout => \ws2812.un1_bit_counter_12_cry_4\,
            clk => \N__27485\,
            ce => 'H',
            sr => \N__27108\
        );

    \ws2812.bit_counter_0_3_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__27855\,
            in1 => \N__24859\,
            in2 => \N__24694\,
            in3 => \N__24682\,
            lcout => \ws2812.bit_counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_4\,
            carryout => \ws2812.un1_bit_counter_12_cry_5\,
            clk => \N__27485\,
            ce => 'H',
            sr => \N__27108\
        );

    \ws2812.bit_counter_2_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24657\,
            in2 => \N__24679\,
            in3 => \N__24637\,
            lcout => \ws2812.bit_counter_6\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_5\,
            carryout => \ws2812.un1_bit_counter_12_cry_6\,
            clk => \N__27485\,
            ce => 'H',
            sr => \N__27108\
        );

    \ws2812.bit_counter_3_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24608\,
            in2 => \N__24634\,
            in3 => \N__24586\,
            lcout => \ws2812.bit_counter_7\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_6\,
            carryout => \ws2812.un1_bit_counter_12_cry_7\,
            clk => \N__27485\,
            ce => 'H',
            sr => \N__27108\
        );

    \ws2812.bit_counter_4_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24834\,
            in2 => \N__24583\,
            in3 => \N__24571\,
            lcout => \ws2812.bit_counter_8\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \ws2812.un1_bit_counter_12_cry_8\,
            clk => \N__27493\,
            ce => 'H',
            sr => \N__27112\
        );

    \ws2812.bit_counter_5_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26354\,
            in2 => \N__24949\,
            in3 => \N__24937\,
            lcout => \ws2812.bit_counter_9\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_8\,
            carryout => \ws2812.un1_bit_counter_12_cry_9\,
            clk => \N__27493\,
            ce => 'H',
            sr => \N__27112\
        );

    \ws2812.bit_counter_0_RNO_0_4_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26403\,
            in2 => \N__24934\,
            in3 => \N__24922\,
            lcout => \ws2812.bit_counter_0_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \ws2812.un1_bit_counter_12_cry_9\,
            carryout => \ws2812.un1_bit_counter_12_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_5_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101011101010"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__24919\,
            in2 => \N__27865\,
            in3 => \N__24910\,
            lcout => \ws2812.bit_counter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27493\,
            ce => 'H',
            sr => \N__27112\
        );

    \ws2812.bit_counter_0_RNIOCUQ_2_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24893\,
            in1 => \N__24832\,
            in2 => \N__26364\,
            in3 => \N__24863\,
            lcout => \ws2812.state_ns_0_i_o2_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNISCT2_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24894\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ws2812.bit_counter_0_RNISCT2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNITDT2_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24864\,
            lcout => \ws2812.bit_counter_0_RNITDT2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNIFOHA_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24833\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ws2812.un6_data_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_0_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__26242\,
            in1 => \N__24982\,
            in2 => \N__25906\,
            in3 => \N__26542\,
            lcout => OPEN,
            ltout => \ws2812.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__24804\,
            in1 => \N__25407\,
            in2 => \N__24814\,
            in3 => \N__26296\,
            lcout => led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27498\,
            ce => 'H',
            sr => \N__27123\
        );

    \ws2812.data_RNO_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__26241\,
            in1 => \N__25276\,
            in2 => \N__25905\,
            in3 => \N__24981\,
            lcout => \ws2812.N_135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI2H7O_2_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25039\,
            in1 => \N__24955\,
            in2 => \_gnd_net_\,
            in3 => \N__28114\,
            lcout => \ws2812.rgb_counter_RNI2H7OZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIFI3M_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28115\,
            in1 => \N__25027\,
            in2 => \_gnd_net_\,
            in3 => \N__25135\,
            lcout => \ws2812.rgb_counter_RNIFI3MZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIDG3M_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26587\,
            in1 => \N__25015\,
            in2 => \_gnd_net_\,
            in3 => \N__28117\,
            lcout => OPEN,
            ltout => \ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIUE972_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__28033\,
            in1 => \N__27933\,
            in2 => \N__25003\,
            in3 => \N__25000\,
            lcout => OPEN,
            ltout => \ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIOQ324_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__27934\,
            in1 => \N__24994\,
            in2 => \N__24988\,
            in3 => \N__24973\,
            lcout => OPEN,
            ltout => \ws2812.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI0NBTB_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27994\,
            in2 => \N__24985\,
            in3 => \N__26533\,
            lcout => \ws2812.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI4J7O_2_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25153\,
            in1 => \N__25114\,
            in2 => \_gnd_net_\,
            in3 => \N__28116\,
            lcout => \ws2812.rgb_counter_RNI4J7OZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_out_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24967\,
            lcout => rgb_data_out_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27505\,
            ce => \N__27194\,
            sr => \N__27128\
        );

    \sb_translator_1.rgb_data_out_13_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => rgb_data_out_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_11_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25147\,
            lcout => rgb_data_out_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_4_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25450\,
            lcout => rgb_data_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_9_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25126\,
            lcout => rgb_data_out_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25633\,
            lcout => rgb_data_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_20_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25084\,
            lcout => rgb_data_out_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25105\,
            lcout => rgb_data_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_out_21_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25096\,
            lcout => rgb_data_out_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27508\,
            ce => \N__27191\,
            sr => \N__27131\
        );

    \sb_translator_1.rgb_data_tmp_20_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25624\,
            in1 => \N__25570\,
            in2 => \N__25534\,
            in3 => \N__25485\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27514\,
            ce => \N__25078\,
            sr => \N__27135\
        );

    \sb_translator_1.rgb_data_tmp_5_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__25866\,
            in1 => \N__25764\,
            in2 => \N__25722\,
            in3 => \N__25663\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27516\,
            ce => \N__25441\,
            sr => \N__27137\
        );

    \sb_translator_1.rgb_data_tmp_4_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25622\,
            in1 => \N__25582\,
            in2 => \N__25538\,
            in3 => \N__25486\,
            lcout => \sb_translator_1.rgb_data_tmpZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27516\,
            ce => \N__25441\,
            sr => \N__27137\
        );

    \ws2812.bit_counter_0_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101111000100"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__26872\,
            in2 => \N__27751\,
            in3 => \N__25274\,
            lcout => \ws2812.bit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27479\,
            ce => 'H',
            sr => \N__27099\
        );

    \ws2812.bit_counter_0_RNIK8UQ_5_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25294\,
            in1 => \N__26392\,
            in2 => \N__25230\,
            in3 => \N__25256\,
            lcout => \ws2812.state_ns_0_i_o2_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNICLHA_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25295\,
            lcout => \ws2812.un6_data_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un6_data_cry_0_c_inv_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__26171\,
            in1 => \N__25257\,
            in2 => \_gnd_net_\,
            in3 => \N__26290\,
            lcout => \ws2812.bit_counter_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIVFT2_5_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25226\,
            lcout => \ws2812.un6_data_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_4_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__27829\,
            in1 => \N__27577\,
            in2 => \_gnd_net_\,
            in3 => \N__25204\,
            lcout => \ws2812.bit_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27486\,
            ce => 'H',
            sr => \N__27109\
        );

    \ws2812.bit_counter_0_0_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__27576\,
            in1 => \N__25195\,
            in2 => \_gnd_net_\,
            in3 => \N__27830\,
            lcout => \ws2812.bit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27486\,
            ce => 'H',
            sr => \N__27109\
        );

    \ws2812.un6_data_cry_0_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26289\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \ws2812.un6_data_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_8_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26278\,
            in2 => \_gnd_net_\,
            in3 => \N__26272\,
            lcout => \ws2812.data_RNOZ0Z_8\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_0\,
            carryout => \ws2812.un6_data_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_9_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26269\,
            in2 => \N__26210\,
            in3 => \N__26263\,
            lcout => \ws2812.data_RNOZ0Z_9\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_1\,
            carryout => \ws2812.un6_data_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_10_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26260\,
            in2 => \N__26208\,
            in3 => \N__26254\,
            lcout => \ws2812.data_RNOZ0Z_10\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_2\,
            carryout => \ws2812.un6_data_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un6_data_cry_3_c_RNIKNFB_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26251\,
            in2 => \N__26211\,
            in3 => \N__26230\,
            lcout => \ws2812.un6_data_cry_3_c_RNIKNFBZ0\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_3\,
            carryout => \ws2812.un6_data_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un6_data_cry_4_c_RNIMQGB_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26227\,
            in2 => \N__26209\,
            in3 => \N__25888\,
            lcout => \ws2812.un6_data_cry_4_c_RNIMQGBZ0\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_4\,
            carryout => \ws2812.un6_data_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_3_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__27696\,
            in1 => \N__25885\,
            in2 => \_gnd_net_\,
            in3 => \N__25879\,
            lcout => \ws2812.data_5_iv_0_47_a2_0_a2_0\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_5\,
            carryout => \ws2812.un6_data_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_11_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25876\,
            in2 => \_gnd_net_\,
            in3 => \N__25870\,
            lcout => \ws2812.data_RNOZ0Z_11\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_6\,
            carryout => \ws2812.un6_data_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_12_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26458\,
            in2 => \_gnd_net_\,
            in3 => \N__26452\,
            lcout => \ws2812.data_RNOZ0Z_12\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \ws2812.un6_data_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_13_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26329\,
            in2 => \_gnd_net_\,
            in3 => \N__26449\,
            lcout => \ws2812.data_RNOZ0Z_13\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_8\,
            carryout => \ws2812.un6_data_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_5_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26374\,
            in2 => \_gnd_net_\,
            in3 => \N__26446\,
            lcout => \ws2812.data_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_9\,
            carryout => \ws2812.un6_data_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_6_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26443\,
            in2 => \_gnd_net_\,
            in3 => \N__26434\,
            lcout => \ws2812.data_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \ws2812.un6_data_cry_10\,
            carryout => \ws2812.un6_data_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26431\,
            in1 => \N__26425\,
            in2 => \N__26419\,
            in3 => \N__26410\,
            lcout => \ws2812.data_5_iv_0_47_a2_0_a2_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_0_RNIUET2_4_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \ws2812.un6_data_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.bit_counter_RNIGPHA_5_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26353\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ws2812.un6_data_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__26323\,
            in1 => \N__26317\,
            in2 => \N__26311\,
            in3 => \N__26302\,
            lcout => \ws2812.data_5_iv_0_47_a2_0_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.data_RNO_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__26578\,
            in1 => \N__26569\,
            in2 => \N__26560\,
            in3 => \N__26548\,
            lcout => \ws2812.data_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIVOJT3_1_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__28032\,
            in1 => \N__27931\,
            in2 => \N__26701\,
            in3 => \N__26485\,
            lcout => OPEN,
            ltout => \ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIUIOE7_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__27932\,
            in1 => \N__26668\,
            in2 => \N__26536\,
            in3 => \N__26818\,
            lcout => \ws2812.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_0_RNIN42Q_3_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__26754\,
            in1 => \N__28106\,
            in2 => \N__26527\,
            in3 => \N__26515\,
            lcout => OPEN,
            ltout => \ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIKHAI1_2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28107\,
            in1 => \N__26506\,
            in2 => \N__26497\,
            in3 => \N__26494\,
            lcout => \ws2812.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un1_rgb_counter_cry_0_c_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27936\,
            in2 => \N__27874\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \ws2812.un1_rgb_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28035\,
            in2 => \N__28006\,
            in3 => \N__26479\,
            lcout => \ws2812.rgb_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ws2812.un1_rgb_counter_cry_0\,
            carryout => \ws2812.un1_rgb_counter_cry_1\,
            clk => \N__27509\,
            ce => 'H',
            sr => \N__27132\
        );

    \ws2812.rgb_counter_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28118\,
            in2 => \N__28048\,
            in3 => \N__26476\,
            lcout => \ws2812.rgb_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ws2812.un1_rgb_counter_cry_1\,
            carryout => \ws2812.un1_rgb_counter_cry_2\,
            clk => \N__27509\,
            ce => 'H',
            sr => \N__27132\
        );

    \ws2812.rgb_counter_RNO_0_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27996\,
            in2 => \N__27949\,
            in3 => \N__26461\,
            lcout => \ws2812.rgb_counter_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \ws2812.un1_rgb_counter_cry_2\,
            carryout => \ws2812.un1_rgb_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_0_3_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__27711\,
            in1 => \N__27861\,
            in2 => \N__26755\,
            in3 => \N__26692\,
            lcout => \ws2812.rgb_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27509\,
            ce => 'H',
            sr => \N__27132\
        );

    \ws2812.rgb_counter_0_RNIP62Q_3_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__26689\,
            in1 => \N__26745\,
            in2 => \N__26617\,
            in3 => \N__28108\,
            lcout => OPEN,
            ltout => \ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIOLAI1_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28109\,
            in1 => \N__26683\,
            in2 => \N__26677\,
            in3 => \N__26674\,
            lcout => \ws2812.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_0_RNIR82Q_3_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__26632\,
            in1 => \N__26659\,
            in2 => \N__28122\,
            in3 => \N__26744\,
            lcout => \ws2812.rgb_data_pmux_6_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_out_2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26647\,
            lcout => rgb_data_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27515\,
            ce => \N__27195\,
            sr => \N__27136\
        );

    \sb_translator_1.rgb_data_out_17_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_data_out_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27517\,
            ce => \N__27192\,
            sr => \N__27138\
        );

    \sb_translator_1.rgb_data_out_23_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26608\,
            lcout => rgb_data_out_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27517\,
            ce => \N__27192\,
            sr => \N__27138\
        );

    \sb_translator_1.rgb_data_out_14_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26599\,
            lcout => rgb_data_out_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27517\,
            ce => \N__27192\,
            sr => \N__27138\
        );

    \sb_translator_1.rgb_data_out_22_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26914\,
            lcout => rgb_data_out_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27517\,
            ce => \N__27192\,
            sr => \N__27138\
        );

    \ws2812.state_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__27562\,
            in1 => \N__27679\,
            in2 => \_gnd_net_\,
            in3 => \N__26904\,
            lcout => \ws2812.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27506\,
            ce => 'H',
            sr => \N__27129\
        );

    \ws2812.rgb_counter_0_RNITA2Q_3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__26800\,
            in1 => \N__26749\,
            in2 => \N__26782\,
            in3 => \N__28112\,
            lcout => OPEN,
            ltout => \ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI0UAI1_2_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28113\,
            in1 => \N__26830\,
            in2 => \N__26821\,
            in3 => \N__26761\,
            lcout => \ws2812.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_out_3_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26812\,
            lcout => rgb_data_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27510\,
            ce => \N__27197\,
            sr => \N__27133\
        );

    \sb_translator_1.rgb_data_out_19_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26794\,
            lcout => rgb_data_out_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27510\,
            ce => \N__27197\,
            sr => \N__27133\
        );

    \sb_translator_1.rgb_data_out_7_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26773\,
            lcout => rgb_data_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27510\,
            ce => \N__27197\,
            sr => \N__27133\
        );

    \ws2812.rgb_counter_RNIRMNJ1_3_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26750\,
            in1 => \N__27995\,
            in2 => \N__28132\,
            in3 => \N__28034\,
            lcout => \ws2812.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNISPAI1_2_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__27526\,
            in1 => \N__28110\,
            in2 => \N__26719\,
            in3 => \N__26707\,
            lcout => \ws2812.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNIGEUO_0_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27935\,
            in2 => \_gnd_net_\,
            in3 => \N__28111\,
            lcout => \ws2812.rgb_counter_0_sqmuxa_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI2AOD3_2_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__27858\,
            in1 => \_gnd_net_\,
            in2 => \N__27742\,
            in3 => \N__28123\,
            lcout => \ws2812.rgb_counter_RNI2AOD3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI19OD3_1_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__28039\,
            in1 => \N__27701\,
            in2 => \_gnd_net_\,
            in3 => \N__27857\,
            lcout => \ws2812.rgb_counter_RNI19OD3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.rgb_counter_RNI3BOD3_3_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__27859\,
            in1 => \N__27997\,
            in2 => \N__27743\,
            in3 => \_gnd_net_\,
            lcout => \ws2812.rgb_counter_RNI3BOD3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.un1_rgb_counter_cry_0_c_RNO_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__27700\,
            lcout => \ws2812.un1_rgb_counter_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ws2812.state_RNIELS35_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27860\,
            in1 => \N__27787\,
            in2 => \N__27744\,
            in3 => \N__27588\,
            lcout => \ws2812.state_RNIELS35Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sb_translator_1.rgb_data_out_6_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27535\,
            lcout => rgb_data_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__27518\,
            ce => \N__27196\,
            sr => \N__27139\
        );
end \INTERFACE\;
