// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 4 2021 00:32:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    reset_n_in,
    led_out,
    mosi_in,
    miso_out,
    cs_n_in,
    clk_spi_in);

    input reset_n_in;
    output led_out;
    input mosi_in;
    output miso_out;
    input cs_n_in;
    input clk_spi_in;

    wire N__28196;
    wire N__28195;
    wire N__28194;
    wire N__28187;
    wire N__28186;
    wire N__28185;
    wire N__28178;
    wire N__28177;
    wire N__28176;
    wire N__28169;
    wire N__28168;
    wire N__28167;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28116;
    wire N__28115;
    wire N__28114;
    wire N__28113;
    wire N__28112;
    wire N__28111;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28107;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28088;
    wire N__28083;
    wire N__28078;
    wire N__28073;
    wire N__28068;
    wire N__28065;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28034;
    wire N__28033;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27936;
    wire N__27935;
    wire N__27934;
    wire N__27933;
    wire N__27932;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27917;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27864;
    wire N__27863;
    wire N__27862;
    wire N__27861;
    wire N__27860;
    wire N__27859;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27855;
    wire N__27852;
    wire N__27845;
    wire N__27842;
    wire N__27831;
    wire N__27830;
    wire N__27829;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27814;
    wire N__27809;
    wire N__27806;
    wire N__27801;
    wire N__27796;
    wire N__27787;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27770;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27758;
    wire N__27751;
    wire N__27750;
    wire N__27749;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27741;
    wire N__27738;
    wire N__27737;
    wire N__27736;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27732;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27719;
    wire N__27716;
    wire N__27715;
    wire N__27712;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27701;
    wire N__27700;
    wire N__27697;
    wire N__27696;
    wire N__27693;
    wire N__27680;
    wire N__27679;
    wire N__27676;
    wire N__27661;
    wire N__27658;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27636;
    wire N__27633;
    wire N__27628;
    wire N__27621;
    wire N__27616;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27589;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27577;
    wire N__27576;
    wire N__27575;
    wire N__27574;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27545;
    wire N__27540;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27519;
    wire N__27518;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27512;
    wire N__27511;
    wire N__27510;
    wire N__27509;
    wire N__27508;
    wire N__27507;
    wire N__27506;
    wire N__27505;
    wire N__27504;
    wire N__27503;
    wire N__27502;
    wire N__27501;
    wire N__27500;
    wire N__27499;
    wire N__27498;
    wire N__27497;
    wire N__27496;
    wire N__27495;
    wire N__27494;
    wire N__27493;
    wire N__27492;
    wire N__27491;
    wire N__27490;
    wire N__27489;
    wire N__27488;
    wire N__27487;
    wire N__27486;
    wire N__27485;
    wire N__27484;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27480;
    wire N__27479;
    wire N__27478;
    wire N__27477;
    wire N__27476;
    wire N__27475;
    wire N__27474;
    wire N__27473;
    wire N__27472;
    wire N__27471;
    wire N__27470;
    wire N__27469;
    wire N__27468;
    wire N__27467;
    wire N__27466;
    wire N__27465;
    wire N__27464;
    wire N__27463;
    wire N__27462;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27457;
    wire N__27456;
    wire N__27455;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27447;
    wire N__27446;
    wire N__27445;
    wire N__27444;
    wire N__27443;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27437;
    wire N__27436;
    wire N__27435;
    wire N__27434;
    wire N__27433;
    wire N__27432;
    wire N__27431;
    wire N__27430;
    wire N__27429;
    wire N__27428;
    wire N__27427;
    wire N__27426;
    wire N__27425;
    wire N__27424;
    wire N__27423;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27419;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27207;
    wire N__27206;
    wire N__27201;
    wire N__27198;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27194;
    wire N__27193;
    wire N__27192;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27159;
    wire N__27158;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27150;
    wire N__27143;
    wire N__27140;
    wire N__27139;
    wire N__27138;
    wire N__27137;
    wire N__27136;
    wire N__27135;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27129;
    wire N__27128;
    wire N__27127;
    wire N__27126;
    wire N__27125;
    wire N__27124;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27116;
    wire N__27115;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27109;
    wire N__27108;
    wire N__27107;
    wire N__27104;
    wire N__27103;
    wire N__27102;
    wire N__27101;
    wire N__27100;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27096;
    wire N__27095;
    wire N__27094;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27087;
    wire N__27086;
    wire N__27085;
    wire N__27084;
    wire N__27083;
    wire N__27082;
    wire N__27081;
    wire N__27080;
    wire N__27079;
    wire N__27078;
    wire N__27077;
    wire N__27076;
    wire N__27075;
    wire N__27074;
    wire N__27073;
    wire N__27072;
    wire N__27071;
    wire N__27070;
    wire N__27069;
    wire N__27068;
    wire N__27067;
    wire N__27066;
    wire N__27065;
    wire N__27064;
    wire N__27063;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26904;
    wire N__26901;
    wire N__26900;
    wire N__26899;
    wire N__26898;
    wire N__26897;
    wire N__26896;
    wire N__26895;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26873;
    wire N__26872;
    wire N__26869;
    wire N__26864;
    wire N__26863;
    wire N__26862;
    wire N__26861;
    wire N__26860;
    wire N__26859;
    wire N__26858;
    wire N__26855;
    wire N__26850;
    wire N__26837;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26745;
    wire N__26744;
    wire N__26741;
    wire N__26736;
    wire N__26733;
    wire N__26728;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26403;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26392;
    wire N__26389;
    wire N__26384;
    wire N__26381;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26354;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26241;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26214;
    wire N__26213;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26192;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26174;
    wire N__26173;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26150;
    wire N__26149;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26137;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26124;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26101;
    wire N__26098;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26078;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26066;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26045;
    wire N__26040;
    wire N__26035;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26023;
    wire N__26016;
    wire N__26013;
    wire N__26006;
    wire N__26003;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25969;
    wire N__25964;
    wire N__25957;
    wire N__25952;
    wire N__25951;
    wire N__25950;
    wire N__25949;
    wire N__25946;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25906;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25866;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25859;
    wire N__25856;
    wire N__25855;
    wire N__25854;
    wire N__25853;
    wire N__25852;
    wire N__25851;
    wire N__25850;
    wire N__25849;
    wire N__25848;
    wire N__25845;
    wire N__25838;
    wire N__25837;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25821;
    wire N__25816;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25792;
    wire N__25789;
    wire N__25782;
    wire N__25777;
    wire N__25774;
    wire N__25765;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25744;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25728;
    wire N__25723;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25715;
    wire N__25712;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25682;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25656;
    wire N__25655;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25582;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25574;
    wire N__25571;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25553;
    wire N__25548;
    wire N__25545;
    wire N__25540;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25504;
    wire N__25499;
    wire N__25494;
    wire N__25491;
    wire N__25486;
    wire N__25485;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25460;
    wire N__25457;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25430;
    wire N__25425;
    wire N__25422;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25407;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25398;
    wire N__25397;
    wire N__25396;
    wire N__25395;
    wire N__25394;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25370;
    wire N__25369;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25361;
    wire N__25360;
    wire N__25357;
    wire N__25356;
    wire N__25355;
    wire N__25352;
    wire N__25347;
    wire N__25342;
    wire N__25339;
    wire N__25326;
    wire N__25319;
    wire N__25312;
    wire N__25311;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25296;
    wire N__25295;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25283;
    wire N__25276;
    wire N__25275;
    wire N__25274;
    wire N__25271;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25253;
    wire N__25248;
    wire N__25245;
    wire N__25240;
    wire N__25231;
    wire N__25230;
    wire N__25227;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25182;
    wire N__25181;
    wire N__25180;
    wire N__25177;
    wire N__25170;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24981;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24906;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24894;
    wire N__24893;
    wire N__24890;
    wire N__24889;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24860;
    wire N__24859;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24838;
    wire N__24835;
    wire N__24834;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24821;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24765;
    wire N__24764;
    wire N__24761;
    wire N__24760;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24741;
    wire N__24738;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24657;
    wire N__24656;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24644;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24612;
    wire N__24609;
    wire N__24608;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24593;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24505;
    wire N__24504;
    wire N__24503;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24488;
    wire N__24479;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24458;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24435;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24431;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24412;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24385;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24360;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24349;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24330;
    wire N__24327;
    wire N__24326;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24304;
    wire N__24301;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24264;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24256;
    wire N__24253;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24225;
    wire N__24220;
    wire N__24219;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24152;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24121;
    wire N__24118;
    wire N__24113;
    wire N__24110;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24093;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24085;
    wire N__24082;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23991;
    wire N__23988;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23955;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23930;
    wire N__23923;
    wire N__23922;
    wire N__23919;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23883;
    wire N__23882;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23771;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23725;
    wire N__23722;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23714;
    wire N__23709;
    wire N__23706;
    wire N__23701;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23629;
    wire N__23626;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23588;
    wire N__23583;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23563;
    wire N__23560;
    wire N__23559;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23551;
    wire N__23548;
    wire N__23543;
    wire N__23540;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23487;
    wire N__23482;
    wire N__23481;
    wire N__23480;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23469;
    wire N__23466;
    wire N__23461;
    wire N__23456;
    wire N__23453;
    wire N__23452;
    wire N__23449;
    wire N__23444;
    wire N__23441;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23426;
    wire N__23425;
    wire N__23424;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23412;
    wire N__23409;
    wire N__23408;
    wire N__23405;
    wire N__23400;
    wire N__23397;
    wire N__23392;
    wire N__23387;
    wire N__23384;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23368;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23362;
    wire N__23357;
    wire N__23352;
    wire N__23347;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23335;
    wire N__23332;
    wire N__23327;
    wire N__23324;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23298;
    wire N__23297;
    wire N__23296;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23273;
    wire N__23272;
    wire N__23267;
    wire N__23264;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23243;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23072;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23050;
    wire N__23047;
    wire N__23042;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23023;
    wire N__23020;
    wire N__23011;
    wire N__23010;
    wire N__23009;
    wire N__23008;
    wire N__23005;
    wire N__23000;
    wire N__22999;
    wire N__22998;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22981;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22959;
    wire N__22954;
    wire N__22945;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22817;
    wire N__22812;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22788;
    wire N__22787;
    wire N__22786;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22782;
    wire N__22781;
    wire N__22780;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22760;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22725;
    wire N__22716;
    wire N__22713;
    wire N__22706;
    wire N__22703;
    wire N__22696;
    wire N__22691;
    wire N__22680;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22652;
    wire N__22645;
    wire N__22644;
    wire N__22643;
    wire N__22640;
    wire N__22639;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22624;
    wire N__22619;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22603;
    wire N__22602;
    wire N__22599;
    wire N__22598;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22564;
    wire N__22561;
    wire N__22560;
    wire N__22557;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22507;
    wire N__22506;
    wire N__22503;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22418;
    wire N__22417;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22405;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22401;
    wire N__22396;
    wire N__22393;
    wire N__22382;
    wire N__22377;
    wire N__22374;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22350;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22337;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22307;
    wire N__22306;
    wire N__22305;
    wire N__22296;
    wire N__22287;
    wire N__22284;
    wire N__22275;
    wire N__22272;
    wire N__22263;
    wire N__22260;
    wire N__22259;
    wire N__22254;
    wire N__22249;
    wire N__22244;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22220;
    wire N__22217;
    wire N__22210;
    wire N__22207;
    wire N__22206;
    wire N__22205;
    wire N__22204;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22193;
    wire N__22176;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22152;
    wire N__22151;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22070;
    wire N__22067;
    wire N__22066;
    wire N__22065;
    wire N__22064;
    wire N__22063;
    wire N__22062;
    wire N__22061;
    wire N__22060;
    wire N__22059;
    wire N__22058;
    wire N__22057;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22051;
    wire N__22050;
    wire N__22049;
    wire N__22048;
    wire N__22047;
    wire N__22046;
    wire N__22045;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22018;
    wire N__22017;
    wire N__22016;
    wire N__22015;
    wire N__22014;
    wire N__22013;
    wire N__22010;
    wire N__22009;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21984;
    wire N__21977;
    wire N__21966;
    wire N__21959;
    wire N__21956;
    wire N__21945;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21905;
    wire N__21898;
    wire N__21891;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21871;
    wire N__21866;
    wire N__21861;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21615;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21517;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21399;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21388;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21373;
    wire N__21364;
    wire N__21363;
    wire N__21362;
    wire N__21361;
    wire N__21360;
    wire N__21357;
    wire N__21356;
    wire N__21353;
    wire N__21352;
    wire N__21345;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21318;
    wire N__21313;
    wire N__21312;
    wire N__21311;
    wire N__21310;
    wire N__21307;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21070;
    wire N__21069;
    wire N__21064;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21052;
    wire N__21049;
    wire N__21042;
    wire N__21035;
    wire N__21030;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20994;
    wire N__20991;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20972;
    wire N__20969;
    wire N__20962;
    wire N__20961;
    wire N__20958;
    wire N__20953;
    wire N__20950;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20932;
    wire N__20929;
    wire N__20920;
    wire N__20917;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20905;
    wire N__20904;
    wire N__20903;
    wire N__20900;
    wire N__20895;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20871;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20865;
    wire N__20862;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20837;
    wire N__20832;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20803;
    wire N__20802;
    wire N__20799;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20787;
    wire N__20782;
    wire N__20781;
    wire N__20780;
    wire N__20777;
    wire N__20776;
    wire N__20775;
    wire N__20766;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20754;
    wire N__20751;
    wire N__20746;
    wire N__20743;
    wire N__20742;
    wire N__20741;
    wire N__20738;
    wire N__20733;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20359;
    wire N__20358;
    wire N__20355;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20320;
    wire N__20319;
    wire N__20318;
    wire N__20317;
    wire N__20316;
    wire N__20313;
    wire N__20312;
    wire N__20309;
    wire N__20302;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20283;
    wire N__20280;
    wire N__20275;
    wire N__20274;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20264;
    wire N__20259;
    wire N__20254;
    wire N__20251;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20227;
    wire N__20226;
    wire N__20223;
    wire N__20222;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20212;
    wire N__20209;
    wire N__20204;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19971;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19956;
    wire N__19953;
    wire N__19948;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19930;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19912;
    wire N__19909;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19895;
    wire N__19894;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19848;
    wire N__19845;
    wire N__19844;
    wire N__19841;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19810;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19771;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19757;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19749;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19654;
    wire N__19653;
    wire N__19652;
    wire N__19651;
    wire N__19646;
    wire N__19645;
    wire N__19644;
    wire N__19643;
    wire N__19642;
    wire N__19637;
    wire N__19634;
    wire N__19625;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19595;
    wire N__19592;
    wire N__19587;
    wire N__19584;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19547;
    wire N__19542;
    wire N__19537;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19529;
    wire N__19524;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19205;
    wire N__19202;
    wire N__19197;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19185;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19163;
    wire N__19156;
    wire N__19153;
    wire N__19152;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19148;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19129;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19097;
    wire N__19096;
    wire N__19095;
    wire N__19090;
    wire N__19085;
    wire N__19082;
    wire N__19075;
    wire N__19074;
    wire N__19073;
    wire N__19072;
    wire N__19071;
    wire N__19062;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19050;
    wire N__19045;
    wire N__19042;
    wire N__19041;
    wire N__19038;
    wire N__19037;
    wire N__19036;
    wire N__19035;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19023;
    wire N__19020;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19004;
    wire N__18997;
    wire N__18996;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18967;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18955;
    wire N__18952;
    wire N__18943;
    wire N__18940;
    wire N__18939;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18926;
    wire N__18919;
    wire N__18916;
    wire N__18915;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18899;
    wire N__18892;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18872;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18858;
    wire N__18857;
    wire N__18856;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18835;
    wire N__18832;
    wire N__18831;
    wire N__18830;
    wire N__18829;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18808;
    wire N__18805;
    wire N__18804;
    wire N__18801;
    wire N__18800;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18786;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18774;
    wire N__18769;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18738;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18728;
    wire N__18723;
    wire N__18722;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18703;
    wire N__18700;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18684;
    wire N__18683;
    wire N__18682;
    wire N__18681;
    wire N__18680;
    wire N__18677;
    wire N__18668;
    wire N__18663;
    wire N__18660;
    wire N__18655;
    wire N__18652;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18644;
    wire N__18643;
    wire N__18638;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18626;
    wire N__18621;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18582;
    wire N__18581;
    wire N__18580;
    wire N__18575;
    wire N__18572;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18564;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18546;
    wire N__18541;
    wire N__18532;
    wire N__18531;
    wire N__18530;
    wire N__18523;
    wire N__18522;
    wire N__18521;
    wire N__18518;
    wire N__18513;
    wire N__18512;
    wire N__18511;
    wire N__18510;
    wire N__18509;
    wire N__18508;
    wire N__18507;
    wire N__18506;
    wire N__18505;
    wire N__18504;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18486;
    wire N__18477;
    wire N__18474;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18427;
    wire N__18426;
    wire N__18425;
    wire N__18424;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18405;
    wire N__18404;
    wire N__18403;
    wire N__18402;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18381;
    wire N__18376;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18368;
    wire N__18363;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18343;
    wire N__18342;
    wire N__18341;
    wire N__18336;
    wire N__18333;
    wire N__18328;
    wire N__18325;
    wire N__18324;
    wire N__18323;
    wire N__18322;
    wire N__18317;
    wire N__18312;
    wire N__18307;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18301;
    wire N__18296;
    wire N__18291;
    wire N__18286;
    wire N__18285;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18273;
    wire N__18270;
    wire N__18263;
    wire N__18260;
    wire N__18253;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18246;
    wire N__18239;
    wire N__18234;
    wire N__18229;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18057;
    wire N__18052;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18031;
    wire N__18028;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17997;
    wire N__17994;
    wire N__17993;
    wire N__17990;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17946;
    wire N__17945;
    wire N__17944;
    wire N__17943;
    wire N__17938;
    wire N__17937;
    wire N__17936;
    wire N__17935;
    wire N__17928;
    wire N__17925;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17905;
    wire N__17904;
    wire N__17901;
    wire N__17898;
    wire N__17893;
    wire N__17892;
    wire N__17891;
    wire N__17884;
    wire N__17881;
    wire N__17880;
    wire N__17879;
    wire N__17876;
    wire N__17875;
    wire N__17872;
    wire N__17865;
    wire N__17860;
    wire N__17857;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17843;
    wire N__17836;
    wire N__17833;
    wire N__17832;
    wire N__17831;
    wire N__17826;
    wire N__17823;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17761;
    wire N__17758;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17750;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17720;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17695;
    wire N__17694;
    wire N__17693;
    wire N__17692;
    wire N__17683;
    wire N__17682;
    wire N__17681;
    wire N__17680;
    wire N__17679;
    wire N__17676;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17660;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17644;
    wire N__17643;
    wire N__17642;
    wire N__17641;
    wire N__17636;
    wire N__17631;
    wire N__17630;
    wire N__17629;
    wire N__17624;
    wire N__17623;
    wire N__17622;
    wire N__17617;
    wire N__17614;
    wire N__17609;
    wire N__17606;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17590;
    wire N__17589;
    wire N__17588;
    wire N__17587;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17557;
    wire N__17552;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17529;
    wire N__17528;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17504;
    wire N__17497;
    wire N__17494;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17451;
    wire N__17450;
    wire N__17449;
    wire N__17448;
    wire N__17447;
    wire N__17444;
    wire N__17443;
    wire N__17432;
    wire N__17427;
    wire N__17424;
    wire N__17419;
    wire N__17418;
    wire N__17417;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17406;
    wire N__17403;
    wire N__17402;
    wire N__17399;
    wire N__17388;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17360;
    wire N__17359;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17347;
    wire N__17346;
    wire N__17343;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17300;
    wire N__17293;
    wire N__17292;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17235;
    wire N__17234;
    wire N__17233;
    wire N__17232;
    wire N__17229;
    wire N__17228;
    wire N__17227;
    wire N__17224;
    wire N__17223;
    wire N__17222;
    wire N__17221;
    wire N__17220;
    wire N__17217;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17203;
    wire N__17202;
    wire N__17201;
    wire N__17200;
    wire N__17199;
    wire N__17198;
    wire N__17197;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17180;
    wire N__17179;
    wire N__17178;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17164;
    wire N__17149;
    wire N__17146;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17116;
    wire N__17107;
    wire N__17106;
    wire N__17105;
    wire N__17104;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17096;
    wire N__17095;
    wire N__17094;
    wire N__17093;
    wire N__17092;
    wire N__17091;
    wire N__17090;
    wire N__17083;
    wire N__17068;
    wire N__17051;
    wire N__17050;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17029;
    wire N__17026;
    wire N__17025;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16918;
    wire N__16917;
    wire N__16916;
    wire N__16915;
    wire N__16912;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16862;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16853;
    wire N__16852;
    wire N__16845;
    wire N__16844;
    wire N__16843;
    wire N__16842;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16807;
    wire N__16800;
    wire N__16789;
    wire N__16786;
    wire N__16785;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16743;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16559;
    wire N__16556;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16539;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16324;
    wire N__16323;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16108;
    wire N__16105;
    wire N__16104;
    wire N__16103;
    wire N__16100;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16083;
    wire N__16078;
    wire N__16077;
    wire N__16072;
    wire N__16071;
    wire N__16070;
    wire N__16067;
    wire N__16062;
    wire N__16057;
    wire N__16054;
    wire N__16053;
    wire N__16050;
    wire N__16049;
    wire N__16046;
    wire N__16039;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16027;
    wire N__16024;
    wire N__16023;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15957;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15933;
    wire N__15932;
    wire N__15929;
    wire N__15928;
    wire N__15925;
    wire N__15924;
    wire N__15923;
    wire N__15918;
    wire N__15913;
    wire N__15908;
    wire N__15901;
    wire N__15900;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15893;
    wire N__15888;
    wire N__15879;
    wire N__15874;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15867;
    wire N__15864;
    wire N__15863;
    wire N__15858;
    wire N__15849;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15823;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15815;
    wire N__15810;
    wire N__15809;
    wire N__15804;
    wire N__15801;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15584;
    wire N__15581;
    wire N__15576;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15554;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15376;
    wire N__15371;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15342;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15158;
    wire N__15155;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15129;
    wire N__15128;
    wire N__15125;
    wire N__15124;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14946;
    wire N__14941;
    wire N__14938;
    wire N__14933;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14911;
    wire N__14908;
    wire N__14907;
    wire N__14906;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14722;
    wire N__14717;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14632;
    wire N__14629;
    wire N__14628;
    wire N__14625;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14605;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14593;
    wire N__14590;
    wire N__14589;
    wire N__14586;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14484;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14473;
    wire N__14472;
    wire N__14471;
    wire N__14470;
    wire N__14463;
    wire N__14460;
    wire N__14453;
    wire N__14450;
    wire N__14443;
    wire N__14442;
    wire N__14439;
    wire N__14438;
    wire N__14437;
    wire N__14436;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14364;
    wire N__14363;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14346;
    wire N__14345;
    wire N__14344;
    wire N__14343;
    wire N__14342;
    wire N__14341;
    wire N__14338;
    wire N__14333;
    wire N__14324;
    wire N__14319;
    wire N__14314;
    wire N__14313;
    wire N__14312;
    wire N__14311;
    wire N__14310;
    wire N__14299;
    wire N__14296;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14284;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14233;
    wire N__14232;
    wire N__14229;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14049;
    wire N__14048;
    wire N__14043;
    wire N__14040;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13992;
    wire N__13991;
    wire N__13990;
    wire N__13989;
    wire N__13988;
    wire N__13987;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13947;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13924;
    wire N__13923;
    wire N__13922;
    wire N__13921;
    wire N__13920;
    wire N__13919;
    wire N__13918;
    wire N__13915;
    wire N__13902;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13872;
    wire N__13869;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13848;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13831;
    wire N__13830;
    wire N__13827;
    wire N__13826;
    wire N__13825;
    wire N__13824;
    wire N__13823;
    wire N__13822;
    wire N__13819;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13802;
    wire N__13799;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13791;
    wire N__13790;
    wire N__13789;
    wire N__13788;
    wire N__13781;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13743;
    wire N__13738;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13666;
    wire N__13665;
    wire N__13664;
    wire N__13663;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13638;
    wire N__13635;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13611;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13566;
    wire N__13561;
    wire N__13554;
    wire N__13551;
    wire N__13544;
    wire N__13541;
    wire N__13536;
    wire N__13531;
    wire N__13526;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13492;
    wire N__13491;
    wire N__13488;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13477;
    wire N__13476;
    wire N__13473;
    wire N__13472;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13461;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13440;
    wire N__13437;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13392;
    wire N__13387;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13360;
    wire N__13355;
    wire N__13348;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13296;
    wire N__13293;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13254;
    wire N__13251;
    wire N__13250;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13210;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13198;
    wire N__13195;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13180;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13168;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13156;
    wire N__13153;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13145;
    wire N__13144;
    wire N__13143;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13128;
    wire N__13127;
    wire N__13126;
    wire N__13125;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13098;
    wire N__13095;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13070;
    wire N__13067;
    wire N__13062;
    wire N__13057;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13035;
    wire N__13030;
    wire N__13029;
    wire N__13028;
    wire N__13025;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13011;
    wire N__13010;
    wire N__13009;
    wire N__13008;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12979;
    wire N__12978;
    wire N__12977;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12937;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12915;
    wire N__12910;
    wire N__12909;
    wire N__12908;
    wire N__12907;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12874;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12856;
    wire N__12851;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12824;
    wire N__12821;
    wire N__12816;
    wire N__12811;
    wire N__12808;
    wire N__12801;
    wire N__12796;
    wire N__12789;
    wire N__12784;
    wire N__12783;
    wire N__12780;
    wire N__12779;
    wire N__12778;
    wire N__12777;
    wire N__12776;
    wire N__12775;
    wire N__12772;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12761;
    wire N__12758;
    wire N__12757;
    wire N__12754;
    wire N__12753;
    wire N__12752;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12705;
    wire N__12698;
    wire N__12693;
    wire N__12692;
    wire N__12683;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12665;
    wire N__12660;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12640;
    wire N__12637;
    wire N__12636;
    wire N__12635;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12584;
    wire N__12577;
    wire N__12574;
    wire N__12569;
    wire N__12566;
    wire N__12561;
    wire N__12554;
    wire N__12547;
    wire N__12540;
    wire N__12537;
    wire N__12532;
    wire N__12531;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12513;
    wire N__12512;
    wire N__12509;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12484;
    wire N__12483;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12442;
    wire N__12439;
    wire N__12438;
    wire N__12435;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12415;
    wire N__12414;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12388;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12376;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12364;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12360;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12327;
    wire N__12326;
    wire N__12325;
    wire N__12324;
    wire N__12323;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12283;
    wire N__12278;
    wire N__12277;
    wire N__12270;
    wire N__12269;
    wire N__12268;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12254;
    wire N__12247;
    wire N__12246;
    wire N__12245;
    wire N__12244;
    wire N__12241;
    wire N__12240;
    wire N__12237;
    wire N__12236;
    wire N__12233;
    wire N__12232;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12203;
    wire N__12202;
    wire N__12199;
    wire N__12198;
    wire N__12195;
    wire N__12194;
    wire N__12191;
    wire N__12190;
    wire N__12187;
    wire N__12186;
    wire N__12183;
    wire N__12182;
    wire N__12179;
    wire N__12178;
    wire N__12175;
    wire N__12174;
    wire N__12171;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12147;
    wire N__12146;
    wire N__12129;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12097;
    wire N__12088;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12061;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12004;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11992;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11980;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11968;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11956;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11944;
    wire N__11943;
    wire N__11942;
    wire N__11941;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11928;
    wire N__11925;
    wire N__11918;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11877;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11815;
    wire N__11812;
    wire N__11807;
    wire N__11798;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11680;
    wire N__11677;
    wire N__11672;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11369;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11331;
    wire N__11330;
    wire N__11329;
    wire N__11328;
    wire N__11325;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10920;
    wire N__10919;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10901;
    wire N__10898;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10867;
    wire N__10864;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10831;
    wire N__10830;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10710;
    wire N__10705;
    wire N__10704;
    wire N__10703;
    wire N__10702;
    wire N__10699;
    wire N__10692;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10615;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10560;
    wire N__10559;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10553;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10531;
    wire N__10530;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10492;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10462;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10447;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10252;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10240;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10228;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10216;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10173;
    wire N__10172;
    wire N__10169;
    wire N__10164;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10122;
    wire N__10117;
    wire N__10114;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10102;
    wire N__10099;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net ;
    wire VCCG0;
    wire \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net ;
    wire GNDG0;
    wire \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net ;
    wire \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net ;
    wire \sb_translator_1.cnt_i_0 ;
    wire bfn_1_3_0_;
    wire \sb_translator_1.cnt_i_1 ;
    wire \sb_translator_1.cnt19_cry_0 ;
    wire \sb_translator_1.cnt_RNIOI3OZ0Z_2 ;
    wire \sb_translator_1.cnt19_cry_1 ;
    wire \sb_translator_1.cnt_RNISN4OZ0Z_3 ;
    wire \sb_translator_1.cnt19_cry_2 ;
    wire \sb_translator_1.cnt_RNI0T5OZ0Z_4 ;
    wire \sb_translator_1.cnt19_cry_3 ;
    wire \sb_translator_1.cnt_RNI427OZ0Z_5 ;
    wire \sb_translator_1.cnt19_cry_4 ;
    wire \sb_translator_1.cnt_RNI878OZ0Z_6 ;
    wire \sb_translator_1.cnt19_cry_5 ;
    wire \sb_translator_1.cnt_RNICC9OZ0Z_7 ;
    wire \sb_translator_1.cnt19_cry_6 ;
    wire \sb_translator_1.cnt19_cry_7 ;
    wire \sb_translator_1.cnt_RNIGHAOZ0Z_8 ;
    wire bfn_1_4_0_;
    wire \sb_translator_1.cnt_RNIKMBOZ0Z_9 ;
    wire \sb_translator_1.cnt19_cry_8 ;
    wire \sb_translator_1.cnt_RNI6O3VZ0Z_10 ;
    wire \sb_translator_1.cnt19_cry_9 ;
    wire \sb_translator_1.cnt_RNIO5UPZ0Z_11 ;
    wire \sb_translator_1.cnt19_cry_10 ;
    wire \sb_translator_1.cnt_RNISAVPZ0Z_12 ;
    wire \sb_translator_1.cnt19_cry_11 ;
    wire \sb_translator_1.cnt_RNI0G0QZ0Z_13 ;
    wire \sb_translator_1.cnt19_cry_12 ;
    wire \sb_translator_1.cnt_RNI4L1QZ0Z_14 ;
    wire \sb_translator_1.cnt19_cry_13 ;
    wire \sb_translator_1.cnt_RNI8Q2QZ0Z_15 ;
    wire \sb_translator_1.cnt19_cry_14 ;
    wire \sb_translator_1.cnt19_cry_15 ;
    wire \sb_translator_1.cnt_i_16 ;
    wire bfn_1_5_0_;
    wire \sb_translator_1.cnt19_cry_16 ;
    wire \sb_translator_1.cnt19_cry_18 ;
    wire \sb_translator_1.cnt19_cry_20 ;
    wire \sb_translator_1.cnt19_cry_21 ;
    wire \sb_translator_1.cnt19_cry_22 ;
    wire \sb_translator_1.cnt19_cry_23 ;
    wire \sb_translator_1.cnt19_cry_24 ;
    wire \sb_translator_1.cnt19_cry_25 ;
    wire bfn_1_6_0_;
    wire \sb_translator_1.cnt19_cry_26 ;
    wire \sb_translator_1.cnt19_cry_27 ;
    wire \sb_translator_1.cnt19_cry_28 ;
    wire \sb_translator_1.cnt19_cry_29 ;
    wire \sb_translator_1.cnt19_cry_30 ;
    wire \sb_translator_1.cnt19_cry_31 ;
    wire \sb_translator_1.cnt19_cry_32 ;
    wire \sb_translator_1.cnt19_cry_33 ;
    wire bfn_1_7_0_;
    wire \sb_translator_1.cnt19_cry_34 ;
    wire \sb_translator_1.cnt19_cry_35 ;
    wire \spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4 ;
    wire \spi_slave_1.un3_mosi_data_out_3 ;
    wire \spi_slave_1.un3_mosi_data_out_3_cascade_ ;
    wire \spi_slave_1.bitcnt_rxZ0Z_0 ;
    wire bfn_1_10_0_;
    wire \spi_slave_1.bitcnt_rxZ0Z_1 ;
    wire \spi_slave_1.bitcnt_rx_cry_0 ;
    wire \spi_slave_1.bitcnt_rxZ0Z_2 ;
    wire \spi_slave_1.bitcnt_rx_cry_1 ;
    wire \spi_slave_1.bitcnt_rxZ0Z_3 ;
    wire \spi_slave_1.bitcnt_rx_cry_2 ;
    wire \spi_slave_1.bitcnt_rx_cry_3 ;
    wire \spi_slave_1.bitcnt_rxZ0Z_4 ;
    wire miso_en;
    wire bfn_1_12_0_;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_0 ;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_1 ;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_2 ;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_3 ;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO ;
    wire \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO ;
    wire \spi_slave_1.mosi_data_inZ0Z_23 ;
    wire \spi_slave_1.mosi_data_inZ0Z_18 ;
    wire \spi_slave_1.mosi_data_inZ0Z_19 ;
    wire \spi_slave_1.mosi_data_inZ0Z_20 ;
    wire \spi_slave_1.mosi_data_inZ0Z_21 ;
    wire \spi_slave_1.mosi_data_inZ0Z_22 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_10 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_2 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_3 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_4 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_5 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_6 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_7 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_8 ;
    wire \sb_translator_1.stateZ0Z_5 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_0_cascade_ ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_13 ;
    wire \sb_translator_1.cntZ0Z_13 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_14 ;
    wire \sb_translator_1.cntZ0Z_14 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_15 ;
    wire \sb_translator_1.cntZ0Z_15 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_16 ;
    wire \sb_translator_1.cntZ0Z_16 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_1 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_11 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_12 ;
    wire \sb_translator_1.cnt_RNO_0Z0Z_9 ;
    wire \sb_translator_1.cntZ0Z_9 ;
    wire \sb_translator_1.cntZ0Z_12 ;
    wire \sb_translator_1.instr_tmpZ0Z_18 ;
    wire \sb_translator_1.instr_tmpZ0Z_19 ;
    wire \sb_translator_1.instr_tmpZ0Z_20 ;
    wire \sb_translator_1.instr_tmpZ0Z_21 ;
    wire \sb_translator_1.instr_tmpZ0Z_22 ;
    wire \sb_translator_1.instr_tmpZ0Z_23 ;
    wire miso_data_in_19;
    wire miso_data_in_20;
    wire miso_data_in_21;
    wire miso_data_in_22;
    wire miso_data_in_23;
    wire miso_data_in_8;
    wire \spi_slave_1.clk_pos_i ;
    wire \spi_slave_1.miso_data_outZ0Z_22 ;
    wire \spi_slave_1.miso_data_outZ0Z_21 ;
    wire \spi_slave_1.m81_ns_1_cascade_ ;
    wire \spi_slave_1.miso_data_outZ0Z_5 ;
    wire \spi_slave_1.miso_data_outZ0Z_4 ;
    wire \spi_slave_1.miso_data_outZ0Z_20 ;
    wire \spi_slave_1.miso_data_outZ0Z_19 ;
    wire \spi_slave_1.m60_ns_1_cascade_ ;
    wire clk_spi;
    wire \spi_slave_1.bitcnt_tx10 ;
    wire \spi_slave_1.bitcnt_tx10_cascade_ ;
    wire \spi_slave_1.miso_data_outZ0Z_8 ;
    wire miso_tx;
    wire \spi_slave_1.N_82 ;
    wire \spi_slave_1.miso_RNOZ0Z_17 ;
    wire \spi_slave_1.miso_RNOZ0Z_10 ;
    wire \spi_slave_1.m48_ns_1_cascade_ ;
    wire \spi_slave_1.N_49_0_cascade_ ;
    wire \spi_slave_1.N_25_0_cascade_ ;
    wire \spi_slave_1.miso_data_outZ0Z_23 ;
    wire \spi_slave_1.miso_data_out_0_sqmuxa ;
    wire \spi_slave_1.N_96_mux ;
    wire \spi_slave_1.N_94_mux ;
    wire \spi_slave_1.N_94_mux_cascade_ ;
    wire \spi_slave_1.bitcnt_txZ0Z_3 ;
    wire \spi_slave_1.N_17_0 ;
    wire \spi_slave_1.N_20_0 ;
    wire \spi_slave_1.N_91 ;
    wire miso;
    wire \spi_slave_1.bitcnt_rxe_0_i ;
    wire \sb_translator_1.un1_num_leds_n_1 ;
    wire bfn_4_3_0_;
    wire \sb_translator_1.un1_num_leds_n_2 ;
    wire \sb_translator_1.un1_num_leds_0_cry_1 ;
    wire \sb_translator_1.un1_num_leds_n_3 ;
    wire \sb_translator_1.un1_num_leds_0_cry_2 ;
    wire \sb_translator_1.un1_num_leds_n_4 ;
    wire \sb_translator_1.un1_num_leds_0_cry_3 ;
    wire \sb_translator_1.un1_num_leds_n_5 ;
    wire \sb_translator_1.un1_num_leds_0_cry_4 ;
    wire \sb_translator_1.un1_num_leds_n_6 ;
    wire \sb_translator_1.un1_num_leds_0_cry_5 ;
    wire \sb_translator_1.un1_num_leds_n_7 ;
    wire \sb_translator_1.un1_num_leds_0_cry_6 ;
    wire \sb_translator_1.un1_num_leds_n_8 ;
    wire \sb_translator_1.un1_num_leds_0_cry_7 ;
    wire \sb_translator_1.un1_num_leds_0_cry_8 ;
    wire \sb_translator_1.un1_num_leds_n_9 ;
    wire bfn_4_4_0_;
    wire \sb_translator_1.un1_num_leds_n_10 ;
    wire \sb_translator_1.un1_num_leds_0_cry_9 ;
    wire \sb_translator_1.un1_num_leds_n_11 ;
    wire \sb_translator_1.un1_num_leds_0_cry_10 ;
    wire \sb_translator_1.un1_num_leds_n_12 ;
    wire \sb_translator_1.un1_num_leds_0_cry_11 ;
    wire \sb_translator_1.un1_num_leds_n_13 ;
    wire \sb_translator_1.un1_num_leds_0_cry_12 ;
    wire \sb_translator_1.un1_num_leds_n_14 ;
    wire \sb_translator_1.un1_num_leds_0_cry_13 ;
    wire \sb_translator_1.un1_num_leds_n_15 ;
    wire \sb_translator_1.un1_num_leds_0_cry_14 ;
    wire \sb_translator_1.un1_num_leds_0_cry_15 ;
    wire \sb_translator_1.un1_num_leds_n_16 ;
    wire \spi_slave_1.mosi_data_inZ0Z_1 ;
    wire reset_n;
    wire reset_n_i;
    wire ram_we_3;
    wire ram_we_13;
    wire \sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_ ;
    wire ram_we_5;
    wire ram_we_7;
    wire ram_we_9;
    wire \sb_translator_1.N_1092 ;
    wire \sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_ ;
    wire ram_we_11;
    wire \sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_ ;
    wire mosi_data_out_17;
    wire demux_data_in_86;
    wire demux_data_in_54;
    wire \demux.N_877_cascade_ ;
    wire demux_data_in_70;
    wire demux_data_in_62;
    wire \demux.N_418_i_0_o2Z0Z_6 ;
    wire demux_data_in_83;
    wire demux_data_in_51;
    wire \demux.N_835_cascade_ ;
    wire demux_data_in_59;
    wire demux_data_in_67;
    wire \demux.N_421_i_0_o2Z0Z_6 ;
    wire demux_data_in_63;
    wire demux_data_in_57;
    wire demux_data_in_87;
    wire demux_data_in_79;
    wire demux_data_in_55;
    wire \demux.N_417_i_0_o2Z0Z_6_cascade_ ;
    wire \demux.N_890 ;
    wire demux_data_in_61;
    wire demux_data_in_77;
    wire demux_data_in_85;
    wire demux_data_in_53;
    wire \demux.N_419_i_0_o2Z0Z_6_cascade_ ;
    wire \demux.N_419_i_0_a3Z0Z_1 ;
    wire demux_data_in_60;
    wire demux_data_in_84;
    wire demux_data_in_76;
    wire demux_data_in_52;
    wire \demux.N_420_i_0_o2Z0Z_6_cascade_ ;
    wire \demux.N_420_i_0_a3Z0Z_1 ;
    wire \spi_slave_1.miso_data_outZ0Z_6 ;
    wire \spi_slave_1.miso_data_outZ0Z_1 ;
    wire \spi_slave_1.miso_data_outZ0Z_3 ;
    wire \spi_slave_1.miso_data_outZ0Z_7 ;
    wire miso_data_in_18;
    wire \spi_slave_1.miso_data_outZ0Z_2 ;
    wire \spi_slave_1.miso_data_outZ0Z_18 ;
    wire \spi_slave_1.m72_ns_1 ;
    wire \spi_slave_1.miso_data_outZ0Z_14 ;
    wire \spi_slave_1.miso_data_outZ0Z_13 ;
    wire \spi_slave_1.bitcnt_txZ0Z_2 ;
    wire \spi_slave_1.miso_RNOZ0Z_12_cascade_ ;
    wire \spi_slave_1.bitcnt_txZ0Z_1 ;
    wire \spi_slave_1.m27_ns_1_cascade_ ;
    wire \spi_slave_1.miso_RNOZ0Z_7 ;
    wire \spi_slave_1.N_28_0 ;
    wire \spi_slave_1.mosi_bufferZ0Z_1 ;
    wire cs_n;
    wire mosi;
    wire \spi_slave_1.mosi_bufferZ0Z_0 ;
    wire \spi_slave_1.clkZ0Z_0 ;
    wire \spi_slave_1.clkZ0Z_1 ;
    wire \spi_slave_1.mosi_data_inZ0Z_17 ;
    wire \spi_slave_1.bitcnt_rxe_0_i_g ;
    wire \spi_slave_1.mosi_data_inZ0Z_9 ;
    wire \spi_slave_1.mosi_data_inZ0Z_8 ;
    wire \spi_slave_1.mosi_data_inZ0Z_10 ;
    wire \spi_slave_1.mosi_data_inZ0Z_11 ;
    wire \spi_slave_1.mosi_data_inZ0Z_12 ;
    wire \spi_slave_1.mosi_data_inZ0Z_13 ;
    wire \spi_slave_1.mosi_data_inZ0Z_14 ;
    wire mosi_data_out_8;
    wire \sb_translator_1.cntZ0Z_0 ;
    wire mosi_data_out_9;
    wire \sb_translator_1.cntZ0Z_1 ;
    wire \sb_translator_1.cntZ0Z_2 ;
    wire mosi_data_out_10;
    wire \spi_slave_1.mosi_data_inZ0Z_16 ;
    wire \spi_slave_1.mosi_data_inZ0Z_3 ;
    wire \spi_slave_1.mosi_data_inZ0Z_2 ;
    wire \spi_slave_1.mosi_data_inZ0Z_5 ;
    wire \spi_slave_1.mosi_data_inZ0Z_6 ;
    wire \spi_slave_1.mosi_data_inZ0Z_7 ;
    wire \spi_slave_1.mosi_data_inZ0Z_4 ;
    wire \spi_slave_1.mosi_data_inZ0Z_0 ;
    wire ram_data_in_0;
    wire ram_data_in_1;
    wire ram_data_in_2;
    wire ram_data_in_3;
    wire ram_data_in_4;
    wire \sb_translator_1.instr_tmpZ1Z_5 ;
    wire mosi_data_out_5;
    wire ram_data_in_5;
    wire \sb_translator_1.instr_tmpZ0Z_6 ;
    wire mosi_data_out_6;
    wire ram_data_in_6;
    wire \sb_translator_1.instr_tmpZ0Z_7 ;
    wire mosi_data_out_7;
    wire ram_data_in_7;
    wire ram_we_0;
    wire ram_we_2;
    wire \sb_translator_1.cnt_RNILAHE_1Z0Z_10 ;
    wire ram_we_10;
    wire ram_we_8;
    wire \sb_translator_1.N_1088 ;
    wire ram_we_12;
    wire \sb_translator_1.cnt_RNILAHE_0Z0Z_10 ;
    wire ram_we_4;
    wire \sb_translator_1.cnt_RNIJ7EF_2Z0Z_9 ;
    wire \sb_translator_1.state_RNI9ILJ_0Z0Z_0 ;
    wire ram_we_6;
    wire \sb_translator_1.cnt_RNIJ7EF_1Z0Z_9 ;
    wire \sb_translator_1.state_RNI9ILJZ0Z_0 ;
    wire ram_we_1;
    wire \sb_translator_1.N_1091_cascade_ ;
    wire \sb_translator_1.N_1089_cascade_ ;
    wire \sb_translator_1.N_1091 ;
    wire \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_ ;
    wire demux_data_in_74;
    wire demux_data_in_82;
    wire demux_data_in_50;
    wire \demux.N_422_i_0_o2Z0Z_6_cascade_ ;
    wire demux_data_in_73;
    wire demux_data_in_81;
    wire demux_data_in_49;
    wire \demux.N_423_i_0_o2Z0Z_6_cascade_ ;
    wire \demux.N_423_i_0_a3Z0Z_1 ;
    wire demux_data_in_58;
    wire \demux.N_422_i_0_a3Z0Z_1 ;
    wire demux_data_in_80;
    wire demux_data_in_72;
    wire demux_data_in_48;
    wire \demux.N_424_i_0_o2_6_cascade_ ;
    wire demux_data_in_56;
    wire \demux.N_424_i_0_a3Z0Z_1 ;
    wire \sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9 ;
    wire \sb_translator_1.state_RNIHS98Z0Z_0 ;
    wire \sb_translator_1.state_RNIHS98_0Z0Z_0 ;
    wire \sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9 ;
    wire \sb_translator_1.N_1089 ;
    wire \demux.N_236_cascade_ ;
    wire \demux.N_235_cascade_ ;
    wire \demux.N_424_i_0_a2Z0Z_6 ;
    wire ram_sel_6;
    wire ram_sel_9;
    wire miso_data_in_9;
    wire \spi_slave_1.miso_data_outZ0Z_17 ;
    wire \spi_slave_1.bitcnt_tx_0_sqmuxa ;
    wire miso_data_in_10;
    wire miso_data_in_11;
    wire miso_data_in_12;
    wire miso_data_in_13;
    wire miso_data_in_14;
    wire miso_data_in_15;
    wire miso_data_in_16;
    wire \sb_translator_1.instr_tmpZ0Z_17 ;
    wire miso_data_in_17;
    wire mosi_data_out_11;
    wire \sb_translator_1.cntZ0Z_3 ;
    wire mosi_data_out_13;
    wire \sb_translator_1.cntZ0Z_5 ;
    wire \sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_9 ;
    wire \sb_translator_1.num_ledsZ0Z_11 ;
    wire \sb_translator_1.num_ledsZ0Z_10 ;
    wire \sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_ ;
    wire \sb_translator_1.ram_sel_6_0_0_a2_0_0_7 ;
    wire \sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10 ;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_0 ;
    wire addr_out_0;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_1 ;
    wire addr_out_1;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_2 ;
    wire addr_out_2;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_3 ;
    wire addr_out_3;
    wire addr_out_4;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_5 ;
    wire addr_out_5;
    wire addr_out_6;
    wire addr_out_7;
    wire \sb_translator_1.cnt_RNILAHE_2Z0Z_10 ;
    wire \sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10 ;
    wire \sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10 ;
    wire mosi_data_out_0;
    wire \sb_translator_1.instr_tmpZ1Z_0 ;
    wire mosi_data_out_1;
    wire \sb_translator_1.instr_tmpZ1Z_1 ;
    wire mosi_data_out_2;
    wire \sb_translator_1.instr_tmpZ1Z_2 ;
    wire mosi_data_out_3;
    wire \sb_translator_1.instr_tmpZ1Z_3 ;
    wire mosi_data_out_4;
    wire \sb_translator_1.instr_tmpZ1Z_4 ;
    wire \sb_translator_1.state_RNIKJOCZ0Z_5 ;
    wire \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ;
    wire \sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11 ;
    wire \sb_translator_1.cnt19_cry_18_THRU_CO ;
    wire \sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_ ;
    wire mosi_rx;
    wire \sb_translator_1.state_RNIOH7V9Z0Z_0 ;
    wire \sb_translator_1.N_58 ;
    wire \sb_translator_1.state_RNIEL0N9_0Z0Z_6 ;
    wire \sb_translator_1.cnt_ram_readZ0Z_0 ;
    wire \sb_translator_1.cnt_ram_readZ0Z_1 ;
    wire demux_data_in_42;
    wire \sb_translator_1.cntZ0Z_11 ;
    wire \sb_translator_1.cntZ0Z_10 ;
    wire \sb_translator_1.ram_we_6_0_0_a2_0_6 ;
    wire miso_data_in_2;
    wire mosi_data_out_22;
    wire \sb_translator_1.N_1087 ;
    wire \sb_translator_1.num_leds_1_sqmuxa_cascade_ ;
    wire \sb_translator_1.send_leds_n_1_sqmuxa ;
    wire \sb_translator_1.N_59 ;
    wire miso_data_in_0;
    wire \sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5 ;
    wire \sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ;
    wire \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0 ;
    wire mosi_data_out_18;
    wire mosi_data_out_19;
    wire mosi_data_out_20;
    wire \sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3 ;
    wire \demux.N_238_cascade_ ;
    wire \demux.N_242_cascade_ ;
    wire \demux.N_424_i_0_a2Z0Z_34_cascade_ ;
    wire \demux.N_424_i_0_aZ0Z2 ;
    wire \demux.N_242 ;
    wire \demux.N_916 ;
    wire ram_sel_5;
    wire \demux.N_916_cascade_ ;
    wire ram_sel_1;
    wire \demux.N_239 ;
    wire \demux.N_241 ;
    wire \demux.N_915 ;
    wire ram_sel_12;
    wire \demux.N_915_cascade_ ;
    wire ram_sel_2;
    wire ram_sel_3;
    wire ram_sel_8;
    wire addr_out_8;
    wire \sb_translator_1.state_RNI88IGAZ0Z_0 ;
    wire \sb_translator_1.state_leds_2_sqmuxa ;
    wire \sb_translator_1.state_ledsZ0 ;
    wire \spi_slave_1.miso_data_outZ0Z_9 ;
    wire \spi_slave_1.miso_data_outZ0Z_10 ;
    wire \spi_slave_1.miso_RNOZ0Z_13 ;
    wire \spi_slave_1.miso_data_outZ0Z_12 ;
    wire \spi_slave_1.miso_data_outZ0Z_11 ;
    wire \spi_slave_1.miso_RNOZ0Z_6 ;
    wire \spi_slave_1.miso_data_outZ0Z_16 ;
    wire \spi_slave_1.miso_data_outZ0Z_0 ;
    wire \spi_slave_1.bitcnt_txZ0Z_4 ;
    wire \spi_slave_1.bitcnt_txZ0Z_0 ;
    wire \spi_slave_1.N_58_0_cascade_ ;
    wire \spi_slave_1.miso_data_outZ0Z_15 ;
    wire \spi_slave_1.N_55_0 ;
    wire \spi_slave_1.mosi_data_inZ0Z_15 ;
    wire \spi_slave_1.un3_mosi_data_out_g ;
    wire \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_5 ;
    wire \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_6 ;
    wire \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_7 ;
    wire \sb_translator_1.num_ledsZ0Z_8 ;
    wire \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_ ;
    wire \sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_3 ;
    wire \sb_translator_1.num_ledsZ0Z_4 ;
    wire \sb_translator_1.cnt19 ;
    wire \sb_translator_1.num_ledsZ0Z_2 ;
    wire \sb_translator_1.state56_a_5_44_cascade_ ;
    wire \sb_translator_1.num_ledsZ0Z_1 ;
    wire \sb_translator_1.cnt_ledsZ0Z_0 ;
    wire bfn_7_4_0_;
    wire \sb_translator_1.cnt_ledsZ0Z_1 ;
    wire \sb_translator_1.cnt_leds_cry_0 ;
    wire \sb_translator_1.cnt_ledsZ0Z_2 ;
    wire \sb_translator_1.cnt_leds_cry_1 ;
    wire \sb_translator_1.cnt_ledsZ0Z_3 ;
    wire \sb_translator_1.cnt_leds_cry_2 ;
    wire \sb_translator_1.cnt_ledsZ0Z_4 ;
    wire \sb_translator_1.cnt_leds_cry_3 ;
    wire \sb_translator_1.cnt_ledsZ0Z_5 ;
    wire \sb_translator_1.cnt_leds_cry_4 ;
    wire \sb_translator_1.cnt_ledsZ0Z_6 ;
    wire \sb_translator_1.cnt_leds_cry_5 ;
    wire \sb_translator_1.cnt_ledsZ0Z_7 ;
    wire \sb_translator_1.cnt_leds_cry_6 ;
    wire \sb_translator_1.cnt_leds_cry_7 ;
    wire \sb_translator_1.cnt_ledsZ0Z_8 ;
    wire bfn_7_5_0_;
    wire \sb_translator_1.cnt_leds_cry_8 ;
    wire \sb_translator_1.cnt_ledsZ0Z_10 ;
    wire \sb_translator_1.cnt_leds_cry_9 ;
    wire \sb_translator_1.cnt_ledsZ0Z_11 ;
    wire \sb_translator_1.cnt_leds_cry_10 ;
    wire \sb_translator_1.cnt_leds_cry_11 ;
    wire \sb_translator_1.cnt_leds_cry_12 ;
    wire \sb_translator_1.cnt_leds_cry_13 ;
    wire \sb_translator_1.cnt_leds_cry_14 ;
    wire \sb_translator_1.cnt_leds_cry_15 ;
    wire bfn_7_6_0_;
    wire \sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1 ;
    wire demux_data_in_40;
    wire demux_data_in_88;
    wire \demux.N_424_i_0_a3Z0Z_4 ;
    wire demux_data_in_8;
    wire \demux.N_424_i_0_o2Z0Z_1_cascade_ ;
    wire demux_data_in_0;
    wire \demux.N_424_i_0_aZ0Z3_cascade_ ;
    wire demux_data_in_35;
    wire demux_data_in_107;
    wire demux_data_in_91;
    wire \demux.N_421_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_2;
    wire demux_data_in_106;
    wire demux_data_in_34;
    wire \demux.N_422_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_90;
    wire \demux.N_422_i_0_a3Z0Z_4 ;
    wire demux_data_in_10;
    wire \demux.N_422_i_0_o2Z0Z_1_cascade_ ;
    wire demux_data_in_9;
    wire demux_data_in_89;
    wire \demux.N_423_i_0_a3Z0Z_5_cascade_ ;
    wire demux_data_in_43;
    wire \demux.N_837 ;
    wire \demux.N_424_i_0_a2Z0Z_34 ;
    wire \demux.N_918_cascade_ ;
    wire demux_data_in_105;
    wire \demux.N_424_i_0_a2Z0Z_5_cascade_ ;
    wire demux_data_in_33;
    wire \demux.N_423_i_0_o2Z0Z_0 ;
    wire \demux.N_918 ;
    wire \demux.N_424_i_0_a2Z0Z_7 ;
    wire \demux.N_424_i_0_o2_0_1 ;
    wire \demux.N_236 ;
    wire \demux.N_235 ;
    wire \demux.N_424_i_0_o2_0Z0Z_2 ;
    wire \demux.N_237 ;
    wire \demux.N_424_i_0_o2_0_8Z0Z_1_cascade_ ;
    wire \demux.N_238 ;
    wire \demux.N_917 ;
    wire \demux.N_424_i_0_o2_0_7_cascade_ ;
    wire \demux.N_424_i_0_o2_0_10 ;
    wire \demux.N_424_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_16;
    wire demux_data_in_96;
    wire demux_data_in_64;
    wire \demux.N_424_i_0_o2Z0Z_4_cascade_ ;
    wire \demux.N_424_i_0_o2Z0Z_8 ;
    wire \demux.N_424_i_0_aZ0Z3 ;
    wire \demux.N_424_i_0_o2_9 ;
    wire \demux.N_424_i_0_o2Z0Z_8_cascade_ ;
    wire \demux.N_424_i_0_o2Z0Z_7 ;
    wire demux_data_in_24;
    wire \demux.N_424_i_0_a3Z0Z_7 ;
    wire ram_sel_0;
    wire ram_sel_11;
    wire \demux.N_906_cascade_ ;
    wire ram_sel_4;
    wire \demux.N_424_i_0_o2_0Z0Z_3 ;
    wire demux_data_in_28;
    wire ram_sel_13;
    wire ram_sel_10;
    wire ram_sel_7;
    wire \demux.N_240 ;
    wire demux_data_in_29;
    wire \sb_translator_1.state56_a_5_ac0_1 ;
    wire bfn_8_3_0_;
    wire \sb_translator_1.cnt_leds_RNIJDTTZ0Z_2 ;
    wire \sb_translator_1.state56_a_5_44 ;
    wire \sb_translator_1.state56_a_5_cry_0_c_THRU_CO ;
    wire \sb_translator_1.cnt_leds_RNIBOUEZ0Z_2 ;
    wire \sb_translator_1.cnt_leds_RNIPJTTZ0Z_3 ;
    wire \sb_translator_1.state56_a_5_cry_0 ;
    wire \sb_translator_1.cnt_leds_RNIERUEZ0Z_3 ;
    wire \sb_translator_1.cnt_leds_RNIVPTTZ0Z_4 ;
    wire \sb_translator_1.state56_a_5_cry_1 ;
    wire \sb_translator_1.cnt_leds_RNIHUUEZ0Z_4 ;
    wire \sb_translator_1.cnt_leds_RNI50UTZ0Z_5 ;
    wire \sb_translator_1.state56_a_5_cry_2 ;
    wire \sb_translator_1.cnt_leds_RNIK1VEZ0Z_5 ;
    wire \sb_translator_1.cnt_leds_RNIB6UTZ0Z_6 ;
    wire \sb_translator_1.state56_a_5_cry_3 ;
    wire \sb_translator_1.cnt_leds_RNIHCUTZ0Z_7 ;
    wire \sb_translator_1.cnt_leds_RNIN4VEZ0Z_6 ;
    wire \sb_translator_1.state56_a_5_cry_4 ;
    wire \sb_translator_1.cnt_leds_RNINIUTZ0Z_8 ;
    wire \sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7 ;
    wire \sb_translator_1.state56_a_5_cry_5 ;
    wire \sb_translator_1.state56_a_5_cry_6 ;
    wire \sb_translator_1.num_leds_RNITOUTZ0Z_8 ;
    wire \sb_translator_1.cnt_leds_RNITAVEZ0Z_8 ;
    wire bfn_8_4_0_;
    wire \sb_translator_1.num_leds_RNIH2E91Z0Z_9 ;
    wire \sb_translator_1.num_leds_RNI0EVEZ0Z_8 ;
    wire \sb_translator_1.state56_a_5_cry_7 ;
    wire \sb_translator_1.num_leds_RNICJVN1Z0Z_10 ;
    wire \sb_translator_1.num_leds_RNIHKEQZ0Z_9 ;
    wire \sb_translator_1.state56_a_5_cry_8 ;
    wire \sb_translator_1.num_leds_RNIP02R1Z0Z_11 ;
    wire \sb_translator_1.num_leds_RNIRUGTZ0Z_10 ;
    wire \sb_translator_1.state56_a_5_cry_9 ;
    wire \sb_translator_1.state56_a_5_cry_10 ;
    wire \sb_translator_1.state56_a_5_cry_11 ;
    wire \sb_translator_1.state56_a_5_cry_12 ;
    wire \sb_translator_1.state56_a_5_cry_13 ;
    wire \sb_translator_1.state56_a_5_cry_14 ;
    wire bfn_8_5_0_;
    wire \sb_translator_1.cnt_ledsZ0Z_16 ;
    wire \sb_translator_1.cnt_leds_i_16_cascade_ ;
    wire \sb_translator_1.num_leds_RNIOJBMZ0Z_15 ;
    wire \sb_translator_1.num_leds_RNIU1HTZ0Z_11 ;
    wire \sb_translator_1.cnt_leds_RNIV62R1Z0Z_13 ;
    wire \sb_translator_1.cnt_leds_RNI48HTZ0Z_14 ;
    wire \sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_ ;
    wire \sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15 ;
    wire \sb_translator_1.num_ledsZ0Z_15 ;
    wire \sb_translator_1.cnt_leds_i_16 ;
    wire \sb_translator_1.cnt_ledsZ0Z_15 ;
    wire \sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15 ;
    wire \sb_translator_1.num_ledsZ0Z_12 ;
    wire \sb_translator_1.cnt_ledsZ0Z_13 ;
    wire \sb_translator_1.cnt_leds_RNI15HTZ0Z_13 ;
    wire \sb_translator_1.num_ledsZ0Z_14 ;
    wire \sb_translator_1.num_ledsZ0Z_13 ;
    wire \sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_ ;
    wire \sb_translator_1.cnt_ledsZ0Z_14 ;
    wire \sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14 ;
    wire demux_data_in_66;
    wire demux_data_in_30;
    wire demux_data_in_102;
    wire demux_data_in_32;
    wire demux_data_in_104;
    wire \demux.N_424_i_0_o2_0Z0Z_0 ;
    wire demux_data_in_44;
    wire demux_data_in_22;
    wire \demux.N_418_i_0_o2Z0Z_4 ;
    wire demux_data_in_78;
    wire \demux.N_884_cascade_ ;
    wire demux_data_in_27;
    wire demux_data_in_19;
    wire demux_data_in_99;
    wire demux_data_in_75;
    wire \demux.N_424_i_0_a2Z0Z_0 ;
    wire \demux.N_421_i_0_o2Z0Z_4_cascade_ ;
    wire \demux.N_421_i_0_a3Z0Z_7 ;
    wire demux_data_in_11;
    wire \demux.N_421_i_0_o2Z0Z_8_cascade_ ;
    wire \demux.N_421_i_0_o2Z0Z_2 ;
    wire \demux.N_422_i_0_o2Z0Z_8 ;
    wire \demux.N_422_i_0_o2Z0Z_9 ;
    wire \demux.N_422_i_0_aZ0Z3 ;
    wire \demux.N_422_i_0_o2Z0Z_7 ;
    wire \sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1 ;
    wire mosi_data_out_16;
    wire \sb_translator_1.cntZ0Z_8 ;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_8 ;
    wire \sb_translator_1.cnt_ledsZ0Z_12 ;
    wire \sb_translator_1.cnt_ledsZ0Z_9 ;
    wire \sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9 ;
    wire demux_data_in_26;
    wire \demux.N_422_i_0_a3Z0Z_7 ;
    wire demux_data_in_15;
    wire demux_data_in_25;
    wire demux_data_in_17;
    wire demux_data_in_97;
    wire demux_data_in_65;
    wire \demux.N_423_i_0_o2Z0Z_4_cascade_ ;
    wire \demux.N_423_i_0_a3Z0Z_7 ;
    wire demux_data_in_41;
    wire \demux.N_423_i_0_o2Z0Z_8_cascade_ ;
    wire \demux.N_423_i_0_o2Z0Z_2 ;
    wire demux_data_in_111;
    wire demux_data_in_39;
    wire demux_data_in_95;
    wire \demux.N_417_i_0_o2Z0Z_0_cascade_ ;
    wire \demux.N_417_i_0_o2Z0Z_1 ;
    wire demux_data_in_47;
    wire \demux.N_417_i_0_a3Z0Z_4 ;
    wire demux_data_in_109;
    wire demux_data_in_37;
    wire demux_data_in_93;
    wire \demux.N_419_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_45;
    wire \demux.N_419_i_0_o2Z0Z_2_cascade_ ;
    wire demux_data_in_13;
    wire \demux.N_419_i_0_a3Z0Z_5 ;
    wire demux_data_in_69;
    wire \demux.N_419_i_0_a3Z0Z_7 ;
    wire \demux.N_419_i_0_o2Z0Z_8 ;
    wire \sb_translator_1.state56_a_5_6 ;
    wire \sb_translator_1.state56_a_5_11 ;
    wire \sb_translator_1.state56_a_5_5 ;
    wire \sb_translator_1.state56_a_5_13 ;
    wire \sb_translator_1.state56_a_5_14 ;
    wire \sb_translator_1.N_318_i_i_o2_12_cascade_ ;
    wire \sb_translator_1.state56_17 ;
    wire \sb_translator_1.state_leds_RNIGMAHZ0 ;
    wire \sb_translator_1.N_318_i_i_o2_15_cascade_ ;
    wire \sb_translator_1.N_712_cascade_ ;
    wire \sb_translator_1.num_leds_1_sqmuxa ;
    wire \sb_translator_1.stateZ0Z_7 ;
    wire \sb_translator_1.state56_a_5_2 ;
    wire \sb_translator_1.state56_a_5_7 ;
    wire \sb_translator_1.N_318_i_i_o2_0 ;
    wire \sb_translator_1.state56_a_5_12 ;
    wire \sb_translator_1.N_318_i_i_o2_8 ;
    wire \sb_translator_1.N_729 ;
    wire \sb_translator_1.N_712 ;
    wire \sb_translator_1.stateZ0Z_0 ;
    wire \sb_translator_1.state_RNIOCIR9Z0Z_5 ;
    wire \sb_translator_1.state56_a_5_4 ;
    wire \sb_translator_1.state56_a_5_10 ;
    wire \sb_translator_1.state56_a_5_3 ;
    wire \sb_translator_1.state56_a_5_16 ;
    wire \sb_translator_1.state56_a_5_8 ;
    wire \sb_translator_1.state56_a_5_9 ;
    wire \sb_translator_1.N_318_i_i_o2_11_cascade_ ;
    wire \sb_translator_1.state56_a_5_15 ;
    wire \sb_translator_1.N_318_i_i_o2_14 ;
    wire \sb_translator_1.state_RNII30CZ0Z_0 ;
    wire \sb_translator_1.stateZ0Z_1 ;
    wire mosi_data_out_23;
    wire mosi_data_out_21;
    wire \sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0 ;
    wire mosi_data_out_12;
    wire \sb_translator_1.cntZ0Z_4 ;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_4 ;
    wire mosi_data_out_14;
    wire \sb_translator_1.cntZ0Z_6 ;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_6 ;
    wire \sb_translator_1.stateZ0Z_6 ;
    wire mosi_data_out_15;
    wire \sb_translator_1.cntZ0Z_7 ;
    wire \sb_translator_1.addr_out_RNO_0Z0Z_7 ;
    wire \ws2812.new_data_req_e_1 ;
    wire \ws2812.N_140_cascade_ ;
    wire ws2812_next_led;
    wire \sb_translator_1.rgb_data_tmpZ0Z_0 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_10 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_12 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_18 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_15 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_16 ;
    wire demux_data_in_94;
    wire demux_data_in_110;
    wire \demux.N_418_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_38;
    wire demux_data_in_46;
    wire \demux.N_418_i_0_o2Z0Z_1_cascade_ ;
    wire \demux.N_424_i_0_a2Z0Z_8 ;
    wire demux_data_in_14;
    wire \demux.N_880 ;
    wire demux_data_in_36;
    wire \demux.N_424_i_0_a2Z0Z_4 ;
    wire \demux.N_424_i_0_a2Z0Z_5 ;
    wire demux_data_in_108;
    wire \demux.N_424_i_0_a2Z0Z_11 ;
    wire \demux.N_420_i_0_o2Z0Z_0_cascade_ ;
    wire demux_data_in_92;
    wire \demux.N_424_i_0_a2Z0Z_2 ;
    wire demux_data_in_12;
    wire \demux.N_420_i_0_o2Z0Z_1_cascade_ ;
    wire \demux.N_420_i_0_a3Z0Z_4 ;
    wire demux_data_in_7;
    wire \demux.N_888_cascade_ ;
    wire demux_data_in_6;
    wire \demux.N_874_cascade_ ;
    wire demux_data_in_4;
    wire \demux.N_417_i_0_o2Z0Z_9 ;
    wire \demux.N_888 ;
    wire \demux.N_417_i_0_o2Z0Z_7 ;
    wire miso_data_in_7;
    wire \demux.N_874 ;
    wire \demux.N_418_i_0_o2Z0Z_8 ;
    wire \demux.N_418_i_0_o2Z0Z_9 ;
    wire \demux.N_418_i_0_o2Z0Z_7 ;
    wire miso_data_in_6;
    wire miso_data_in_5;
    wire \demux.N_421_i_0_o2Z0Z_9 ;
    wire demux_data_in_3;
    wire \demux.N_421_i_0_o2Z0Z_10 ;
    wire miso_data_in_3;
    wire \demux.N_423_i_0_o2Z0Z_9 ;
    wire demux_data_in_1;
    wire \demux.N_423_i_0_o2Z0Z_10 ;
    wire miso_data_in_1;
    wire miso_data_in_4;
    wire \sb_translator_1.state_g_1 ;
    wire demux_data_in_31;
    wire \demux.N_424_i_0_a2Z0Z_1 ;
    wire demux_data_in_71;
    wire \demux.N_417_i_0_a3Z0Z_7_cascade_ ;
    wire \demux.N_417_i_0_o2Z0Z_8 ;
    wire demux_data_in_103;
    wire demux_data_in_23;
    wire \demux.N_417_i_0_o2Z0Z_4 ;
    wire demux_data_in_18;
    wire demux_data_in_98;
    wire \demux.N_422_i_0_o2Z0Z_4 ;
    wire demux_data_in_101;
    wire demux_data_in_21;
    wire \demux.N_419_i_0_o2Z0Z_4 ;
    wire demux_data_in_100;
    wire \demux.N_424_i_0_a2Z0Z_3 ;
    wire demux_data_in_20;
    wire \demux.N_424_i_0_a2Z0Z_10 ;
    wire demux_data_in_68;
    wire \demux.N_424_i_0_a2Z0Z_9 ;
    wire \demux.N_420_i_0_o2Z0Z_4_cascade_ ;
    wire \demux.N_420_i_0_a3Z0Z_7 ;
    wire \ws2812.state_ns_0_i_o2_6_0_cascade_ ;
    wire \ws2812.N_105_cascade_ ;
    wire \ws2812.state_ns_0_i_o2_6_0 ;
    wire \ws2812.un1_bit_counter_12_cry_0_c_RNOZ0 ;
    wire bfn_11_5_0_;
    wire \ws2812.bit_counter_RNI5NQB3Z0Z_1 ;
    wire \ws2812.un1_bit_counter_12_cry_0 ;
    wire \ws2812.bit_counter_0_RNIJC643Z0Z_0 ;
    wire \ws2812.un1_bit_counter_12_cry_1 ;
    wire \ws2812.bit_counterZ0Z_3 ;
    wire \ws2812.bit_counter_0_RNIKD643Z0Z_1 ;
    wire \ws2812.bit_counter_0_RNO_0Z0Z_1 ;
    wire \ws2812.un1_bit_counter_12_cry_2 ;
    wire \ws2812.bit_counter_0_RNILE643Z0Z_2 ;
    wire \ws2812.un1_bit_counter_12_cry_3 ;
    wire \ws2812.bit_counter_0_RNIMF643Z0Z_3 ;
    wire \ws2812.un1_bit_counter_12_cry_4 ;
    wire \ws2812.bit_counter_RNI6OQB3Z0Z_2 ;
    wire \ws2812.bit_counter_6 ;
    wire \ws2812.un1_bit_counter_12_cry_5 ;
    wire \ws2812.bit_counter_RNI7PQB3Z0Z_3 ;
    wire \ws2812.bit_counter_7 ;
    wire \ws2812.un1_bit_counter_12_cry_6 ;
    wire \ws2812.un1_bit_counter_12_cry_7 ;
    wire \ws2812.bit_counter_RNI8QQB3Z0Z_4 ;
    wire bfn_11_6_0_;
    wire \ws2812.bit_counter_RNI9RQB3Z0Z_5 ;
    wire \ws2812.un1_bit_counter_12_cry_8 ;
    wire \ws2812.bit_counter_0_RNING643Z0Z_4 ;
    wire \ws2812.un1_bit_counter_12_cry_9 ;
    wire \ws2812.un1_bit_counter_12_axb_11 ;
    wire \ws2812.un1_bit_counter_12_cry_10 ;
    wire \ws2812.state_ns_0_i_o2_7_0 ;
    wire \ws2812.bit_counterZ0Z_4 ;
    wire \ws2812.bit_counterZ0Z_5 ;
    wire \ws2812.bit_counter_8 ;
    wire \ws2812.N_52_cascade_ ;
    wire led;
    wire rgb_data_out_12;
    wire rgb_data_out_15;
    wire rgb_data_out_10;
    wire \ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_ ;
    wire \ws2812.rgb_counter_RNI2H7OZ0Z_2 ;
    wire \ws2812.rgb_counter_RNIFI3MZ0Z_2 ;
    wire \ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_ ;
    wire \ws2812.N_108_cascade_ ;
    wire \ws2812.N_107 ;
    wire \ws2812.rgb_counter_RNI4J7OZ0Z_2 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_8 ;
    wire rgb_data_out_8;
    wire \sb_translator_1.rgb_data_tmpZ0Z_13 ;
    wire rgb_data_out_13;
    wire \sb_translator_1.rgb_data_tmpZ0Z_11 ;
    wire rgb_data_out_11;
    wire \sb_translator_1.rgb_data_tmpZ0Z_9 ;
    wire rgb_data_out_9;
    wire \sb_translator_1.rgb_data_tmpZ0Z_1 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_21 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_20 ;
    wire \sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1 ;
    wire \demux.N_424_i_0_o2Z0Z_0 ;
    wire \demux.N_419_i_0_o2Z0Z_9 ;
    wire demux_data_in_5;
    wire \demux.N_419_i_0_o2Z0Z_10 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_5 ;
    wire \demux.N_420_i_0_o2Z0Z_8 ;
    wire \demux.N_420_i_0_o2Z0Z_9 ;
    wire \demux.N_420_i_0_aZ0Z3 ;
    wire \demux.N_420_i_0_o2Z0Z_7 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_4 ;
    wire \sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1 ;
    wire \ws2812.stateZ0Z_1 ;
    wire \ws2812.state_ns_0_i_o2_8_0 ;
    wire \ws2812.bit_counterZ0Z_1 ;
    wire \ws2812.bit_counterZ0Z_0 ;
    wire \ws2812.bit_counter_11 ;
    wire \ws2812.bit_counter_0_RNO_0Z0Z_4 ;
    wire \ws2812.bit_counter_0_RNO_0Z0Z_0 ;
    wire \ws2812.bit_counterZ0Z_2 ;
    wire \ws2812.bit_counter_i_0 ;
    wire bfn_12_5_0_;
    wire \ws2812.un6_data_axb_1 ;
    wire \ws2812.un6_data_cry_0 ;
    wire \ws2812.bit_counter_0_RNIQAT2Z0Z_0 ;
    wire \ws2812.un6_data_cry_1 ;
    wire \ws2812.bit_counter_0_RNIRBT2Z0Z_1 ;
    wire \ws2812.un6_data_cry_2 ;
    wire \ws2812.bit_counter_0_RNISCT2Z0Z_2 ;
    wire \ws2812.un6_data_cry_3_c_RNIKNFBZ0 ;
    wire \ws2812.un6_data_cry_3 ;
    wire \ws2812.bit_counter_0_RNITDT2Z0Z_3 ;
    wire CONSTANT_ONE_NET;
    wire \ws2812.un6_data_cry_4_c_RNIMQGBZ0 ;
    wire \ws2812.un6_data_cry_4 ;
    wire \ws2812.un6_data_axb_6 ;
    wire \ws2812.un6_data_cry_5 ;
    wire \ws2812.un6_data_axb_7 ;
    wire \ws2812.un6_data_cry_6 ;
    wire \ws2812.un6_data_cry_7 ;
    wire \ws2812.un6_data_axb_8 ;
    wire bfn_12_6_0_;
    wire \ws2812.un6_data_cry_8 ;
    wire \ws2812.un6_data_cry_9 ;
    wire \ws2812.un6_data_axb_11 ;
    wire \ws2812.un6_data_cry_10 ;
    wire \ws2812.data_RNOZ0Z_11 ;
    wire \ws2812.data_RNOZ0Z_12 ;
    wire \ws2812.data_RNOZ0Z_13 ;
    wire \ws2812.un6_data_cry_11 ;
    wire \ws2812.bit_counter_10 ;
    wire \ws2812.un6_data_axb_10 ;
    wire \ws2812.bit_counter_9 ;
    wire \ws2812.un6_data_axb_9 ;
    wire \ws2812.data_RNOZ0Z_6 ;
    wire \ws2812.data_RNOZ0Z_5 ;
    wire \ws2812.data_5_iv_0_47_a2_0_a2_0 ;
    wire \ws2812.data_5_iv_0_47_a2_0_a2_6_1 ;
    wire \ws2812.data_5_iv_0_47_a2_0_a2_6 ;
    wire \ws2812.data_RNOZ0Z_10 ;
    wire \ws2812.data_RNOZ0Z_9 ;
    wire \ws2812.data_RNOZ0Z_8 ;
    wire \ws2812.N_135 ;
    wire \ws2812.data_RNOZ0Z_2 ;
    wire \ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_ ;
    wire \ws2812.N_115 ;
    wire rgb_data_out_16;
    wire rgb_data_out_0;
    wire rgb_data_out_20;
    wire \ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_ ;
    wire rgb_data_out_4;
    wire \ws2812.N_127 ;
    wire bfn_12_8_0_;
    wire \ws2812.un1_rgb_counter_cry_0 ;
    wire \ws2812.un1_rgb_counter_cry_1 ;
    wire \ws2812.rgb_counter_RNO_0Z0Z_3 ;
    wire \ws2812.un1_rgb_counter_cry_2 ;
    wire \ws2812.un1_rgb_counter_cry_3 ;
    wire rgb_data_out_1;
    wire rgb_data_out_21;
    wire \ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_ ;
    wire rgb_data_out_5;
    wire \ws2812.N_120 ;
    wire rgb_data_out_18;
    wire \sb_translator_1.rgb_data_tmpZ0Z_2 ;
    wire rgb_data_out_2;
    wire \sb_translator_1.rgb_data_tmpZ0Z_17 ;
    wire rgb_data_out_17;
    wire \sb_translator_1.rgb_data_tmpZ0Z_23 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_14 ;
    wire rgb_data_out_14;
    wire \sb_translator_1.rgb_data_tmpZ0Z_22 ;
    wire \ws2812.N_105 ;
    wire rgb_data_out_23;
    wire \ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_ ;
    wire \ws2812.N_117 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_3 ;
    wire rgb_data_out_3;
    wire \sb_translator_1.rgb_data_tmpZ0Z_19 ;
    wire rgb_data_out_19;
    wire \sb_translator_1.rgb_data_tmpZ0Z_7 ;
    wire rgb_data_out_7;
    wire \ws2812.rgb_counter_4 ;
    wire rgb_data_out_22;
    wire \ws2812.rgb_data_pmux_6_i_m2_ns_1 ;
    wire \ws2812.N_124 ;
    wire \ws2812.rgb_counter_0_sqmuxa_0_a2_0_1 ;
    wire \ws2812.rgb_counterZ0Z_2 ;
    wire \ws2812.rgb_counter_RNI2AOD3Z0Z_2 ;
    wire \ws2812.rgb_counterZ0Z_1 ;
    wire \ws2812.rgb_counter_RNI19OD3Z0Z_1 ;
    wire \ws2812.rgb_counterZ0Z_3 ;
    wire \ws2812.rgb_counter_RNI3BOD3Z0Z_3 ;
    wire \ws2812.rgb_counterZ0Z_0 ;
    wire \ws2812.un1_rgb_counter_cry_0_c_RNOZ0 ;
    wire \ws2812.N_106 ;
    wire send_leds_n;
    wire \ws2812.stateZ0Z_0 ;
    wire \ws2812.N_228 ;
    wire \ws2812.state_RNIELS35Z0Z_0 ;
    wire \sb_translator_1.rgb_data_tmpZ0Z_6 ;
    wire rgb_data_out_6;
    wire _gnd_net_;
    wire clk_sb;
    wire \sb_translator_1.state_leds_2_sqmuxa_g ;
    wire reset_n_i_g;

    defparam \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_1__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,demux_data_in_15,dangling_wire_1,demux_data_in_14,dangling_wire_2,demux_data_in_13,dangling_wire_3,demux_data_in_12,dangling_wire_4,demux_data_in_11,dangling_wire_5,demux_data_in_10,dangling_wire_6,demux_data_in_9,dangling_wire_7,demux_data_in_8}),
            .RADDR({dangling_wire_8,dangling_wire_9,N__18112,N__16216,N__16432,N__16633,N__14785,N__15004,N__15232,N__15451,N__15655}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__18115,N__16210,N__16426,N__16660,N__14788,N__15013,N__15259,N__15454,N__15688}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,N__13492,dangling_wire_29,N__13671,dangling_wire_30,N__13818,dangling_wire_31,N__12641,dangling_wire_32,N__12753,dangling_wire_33,N__12909,dangling_wire_34,N__13028,dangling_wire_35,N__13143}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26207),
            .WCLKE(N__13897),
            .WCLK(N__27513),
            .WE(N__26214));
    defparam \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_2__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_36,demux_data_in_23,dangling_wire_37,demux_data_in_22,dangling_wire_38,demux_data_in_21,dangling_wire_39,demux_data_in_20,dangling_wire_40,demux_data_in_19,dangling_wire_41,demux_data_in_18,dangling_wire_42,demux_data_in_17,dangling_wire_43,demux_data_in_16}),
            .RADDR({dangling_wire_44,dangling_wire_45,N__18088,N__16192,N__16408,N__16609,N__14760,N__14980,N__15208,N__15427,N__15631}),
            .WADDR({dangling_wire_46,dangling_wire_47,N__18091,N__16186,N__16402,N__16636,N__14763,N__14989,N__15235,N__15430,N__15664}),
            .MASK({dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63}),
            .WDATA({dangling_wire_64,N__13471,dangling_wire_65,N__13672,dangling_wire_66,N__13830,dangling_wire_67,N__12653,dangling_wire_68,N__12776,dangling_wire_69,N__12910,dangling_wire_70,N__13029,dangling_wire_71,N__13144}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26212),
            .WCLKE(N__13324),
            .WCLK(N__27520),
            .WE(N__26218));
    defparam \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_10__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_72,demux_data_in_87,dangling_wire_73,demux_data_in_86,dangling_wire_74,demux_data_in_85,dangling_wire_75,demux_data_in_84,dangling_wire_76,demux_data_in_83,dangling_wire_77,demux_data_in_82,dangling_wire_78,demux_data_in_81,dangling_wire_79,demux_data_in_80}),
            .RADDR({dangling_wire_80,dangling_wire_81,N__18208,N__16310,N__16526,N__16727,N__14881,N__15100,N__15326,N__15547,N__15751}),
            .WADDR({dangling_wire_82,dangling_wire_83,N__18211,N__16306,N__16522,N__16744,N__14884,N__15109,N__15343,N__15550,N__15777}),
            .MASK({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99}),
            .WDATA({dangling_wire_100,N__13491,dangling_wire_101,N__13670,dangling_wire_102,N__13798,dangling_wire_103,N__12654,dangling_wire_104,N__12757,dangling_wire_105,N__12906,dangling_wire_106,N__13024,dangling_wire_107,N__13152}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26156),
            .WCLKE(N__13288),
            .WCLK(N__27463),
            .WE(N__26170));
    defparam \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_5__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_108,demux_data_in_47,dangling_wire_109,demux_data_in_46,dangling_wire_110,demux_data_in_45,dangling_wire_111,demux_data_in_44,dangling_wire_112,demux_data_in_43,dangling_wire_113,demux_data_in_42,dangling_wire_114,demux_data_in_41,dangling_wire_115,demux_data_in_40}),
            .RADDR({dangling_wire_116,dangling_wire_117,N__18178,N__16261,N__16477,N__16678,N__14863,N__15091,N__15277,N__15505,N__15718}),
            .WADDR({dangling_wire_118,dangling_wire_119,N__18181,N__16279,N__16495,N__16699,N__14878,N__15082,N__15298,N__15508,N__15745}),
            .MASK({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .WDATA({dangling_wire_136,N__13440,dangling_wire_137,N__13611,dangling_wire_138,N__13788,dangling_wire_139,N__12635,dangling_wire_140,N__12692,dangling_wire_141,N__12856,dangling_wire_142,N__12948,dangling_wire_143,N__13070}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26066),
            .WCLKE(N__11197),
            .WCLK(N__27431),
            .WE(N__26125));
    defparam \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_11__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_144,demux_data_in_95,dangling_wire_145,demux_data_in_94,dangling_wire_146,demux_data_in_93,dangling_wire_147,demux_data_in_92,dangling_wire_148,demux_data_in_91,dangling_wire_149,demux_data_in_90,dangling_wire_150,demux_data_in_89,dangling_wire_151,demux_data_in_88}),
            .RADDR({dangling_wire_152,dangling_wire_153,N__18184,N__16288,N__16504,N__16705,N__14857,N__15076,N__15304,N__15523,N__15727}),
            .WADDR({dangling_wire_154,dangling_wire_155,N__18187,N__16282,N__16498,N__16730,N__14860,N__15085,N__15329,N__15526,N__15760}),
            .MASK({dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171}),
            .WDATA({dangling_wire_172,N__13472,dangling_wire_173,N__13645,dangling_wire_174,N__13789,dangling_wire_175,N__12642,dangling_wire_176,N__12775,dangling_wire_177,N__12907,dangling_wire_178,N__12977,dangling_wire_179,N__13098}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26172),
            .WCLKE(N__11353),
            .WCLK(N__27478),
            .WE(N__26196));
    defparam \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_0__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_180,demux_data_in_7,dangling_wire_181,demux_data_in_6,dangling_wire_182,demux_data_in_5,dangling_wire_183,demux_data_in_4,dangling_wire_184,demux_data_in_3,dangling_wire_185,demux_data_in_2,dangling_wire_186,demux_data_in_1,dangling_wire_187,demux_data_in_0}),
            .RADDR({dangling_wire_188,dangling_wire_189,N__18228,N__16324,N__16540,N__16743,N__14905,N__15124,N__15342,N__15561,N__15773}),
            .WADDR({dangling_wire_190,dangling_wire_191,N__18229,N__16323,N__16539,N__16750,N__14906,N__15129,N__15349,N__15562,N__15784}),
            .MASK({dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207}),
            .WDATA({dangling_wire_208,N__13487,dangling_wire_209,N__13669,dangling_wire_210,N__13822,dangling_wire_211,N__12655,dangling_wire_212,N__12777,dangling_wire_213,N__12896,dangling_wire_214,N__13030,dangling_wire_215,N__13156}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26155),
            .WCLKE(N__13339),
            .WCLK(N__27447),
            .WE(N__26097));
    defparam \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_4__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_216,demux_data_in_39,dangling_wire_217,demux_data_in_38,dangling_wire_218,demux_data_in_37,dangling_wire_219,demux_data_in_36,dangling_wire_220,demux_data_in_35,dangling_wire_221,demux_data_in_34,dangling_wire_222,demux_data_in_33,dangling_wire_223,demux_data_in_32}),
            .RADDR({dangling_wire_224,dangling_wire_225,N__18202,N__16285,N__16501,N__16702,N__14887,N__15115,N__15301,N__15529,N__15742}),
            .WADDR({dangling_wire_226,dangling_wire_227,N__18205,N__16303,N__16519,N__16723,N__14902,N__15106,N__15322,N__15532,N__15767}),
            .MASK({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243}),
            .WDATA({dangling_wire_244,N__13460,dangling_wire_245,N__13634,dangling_wire_246,N__13823,dangling_wire_247,N__12636,dangling_wire_248,N__12771,dangling_wire_249,N__12873,dangling_wire_250,N__12986,dangling_wire_251,N__13107}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__25951),
            .WCLKE(N__14035),
            .WCLK(N__27424),
            .WE(N__26034));
    defparam \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_6__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_252,demux_data_in_55,dangling_wire_253,demux_data_in_54,dangling_wire_254,demux_data_in_53,dangling_wire_255,demux_data_in_52,dangling_wire_256,demux_data_in_51,dangling_wire_257,demux_data_in_50,dangling_wire_258,demux_data_in_49,dangling_wire_259,demux_data_in_48}),
            .RADDR({dangling_wire_260,dangling_wire_261,N__18154,N__16237,N__16453,N__16654,N__14839,N__15067,N__15253,N__15481,N__15694}),
            .WADDR({dangling_wire_262,dangling_wire_263,N__18157,N__16255,N__16471,N__16675,N__14854,N__15058,N__15274,N__15484,N__15721}),
            .MASK({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279}),
            .WDATA({dangling_wire_280,N__13450,dangling_wire_281,N__13624,dangling_wire_282,N__13802,dangling_wire_283,N__12630,dangling_wire_284,N__12761,dangling_wire_285,N__12866,dangling_wire_286,N__12978,dangling_wire_287,N__13099}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26177),
            .WCLKE(N__13969),
            .WCLK(N__27443),
            .WE(N__26078));
    defparam \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_3__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_288,demux_data_in_31,dangling_wire_289,demux_data_in_30,dangling_wire_290,demux_data_in_29,dangling_wire_291,demux_data_in_28,dangling_wire_292,demux_data_in_27,dangling_wire_293,demux_data_in_26,dangling_wire_294,demux_data_in_25,dangling_wire_295,demux_data_in_24}),
            .RADDR({dangling_wire_296,dangling_wire_297,N__18226,N__16309,N__16525,N__16726,N__14907,N__15130,N__15325,N__15553,N__15766}),
            .WADDR({dangling_wire_298,dangling_wire_299,N__18227,N__16322,N__16538,N__16742,N__14911,N__15128,N__15341,N__15554,N__15780}),
            .MASK({dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .WDATA({dangling_wire_316,N__13484,dangling_wire_317,N__13662,dangling_wire_318,N__13824,dangling_wire_319,N__12652,dangling_wire_320,N__12783,dangling_wire_321,N__12897,dangling_wire_322,N__13009,dangling_wire_323,N__13127}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__25949),
            .WCLKE(N__11230),
            .WCLK(N__27420),
            .WE(N__25950));
    defparam \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_13__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_324,demux_data_in_111,dangling_wire_325,demux_data_in_110,dangling_wire_326,demux_data_in_109,dangling_wire_327,demux_data_in_108,dangling_wire_328,demux_data_in_107,dangling_wire_329,demux_data_in_106,dangling_wire_330,demux_data_in_105,dangling_wire_331,demux_data_in_104}),
            .RADDR({dangling_wire_332,dangling_wire_333,N__18136,N__16240,N__16456,N__16657,N__14809,N__15028,N__15256,N__15475,N__15679}),
            .WADDR({dangling_wire_334,dangling_wire_335,N__18139,N__16234,N__16450,N__16684,N__14812,N__15037,N__15283,N__15478,N__15712}),
            .MASK({dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .WDATA({dangling_wire_352,N__13476,dangling_wire_353,N__13665,dangling_wire_354,N__13791,dangling_wire_355,N__12640,dangling_wire_356,N__12752,dangling_wire_357,N__12905,dangling_wire_358,N__13011,dangling_wire_359,N__13145}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26191),
            .WCLKE(N__11215),
            .WCLK(N__27503),
            .WE(N__26213));
    defparam \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_12__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_360,demux_data_in_103,dangling_wire_361,demux_data_in_102,dangling_wire_362,demux_data_in_101,dangling_wire_363,demux_data_in_100,dangling_wire_364,demux_data_in_99,dangling_wire_365,demux_data_in_98,dangling_wire_366,demux_data_in_97,dangling_wire_367,demux_data_in_96}),
            .RADDR({dangling_wire_368,dangling_wire_369,N__18160,N__16264,N__16480,N__16681,N__14833,N__15052,N__15280,N__15499,N__15703}),
            .WADDR({dangling_wire_370,dangling_wire_371,N__18163,N__16258,N__16474,N__16708,N__14836,N__15061,N__15307,N__15502,N__15736}),
            .MASK({dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387}),
            .WDATA({dangling_wire_388,N__13477,dangling_wire_389,N__13655,dangling_wire_390,N__13790,dangling_wire_391,N__12643,dangling_wire_392,N__12751,dangling_wire_393,N__12904,dangling_wire_394,N__13010,dangling_wire_395,N__13128}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26173),
            .WCLKE(N__13237),
            .WCLK(N__27492),
            .WE(N__26197));
    defparam \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_7__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_396,demux_data_in_63,dangling_wire_397,demux_data_in_62,dangling_wire_398,demux_data_in_61,dangling_wire_399,demux_data_in_60,dangling_wire_400,demux_data_in_59,dangling_wire_401,demux_data_in_58,dangling_wire_402,demux_data_in_57,dangling_wire_403,demux_data_in_56}),
            .RADDR({dangling_wire_404,dangling_wire_405,N__18130,N__16213,N__16429,N__16630,N__14815,N__15043,N__15229,N__15457,N__15670}),
            .WADDR({dangling_wire_406,dangling_wire_407,N__18133,N__16231,N__16447,N__16651,N__14830,N__15034,N__15250,N__15460,N__15697}),
            .MASK({dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423}),
            .WDATA({dangling_wire_424,N__13464,dangling_wire_425,N__13638,dangling_wire_426,N__13825,dangling_wire_427,N__12631,dangling_wire_428,N__12778,dangling_wire_429,N__12895,dangling_wire_430,N__12979,dangling_wire_431,N__13100}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26178),
            .WCLKE(N__11191),
            .WCLK(N__27455),
            .WE(N__26148));
    defparam \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_8__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_432,demux_data_in_71,dangling_wire_433,demux_data_in_70,dangling_wire_434,demux_data_in_69,dangling_wire_435,demux_data_in_68,dangling_wire_436,demux_data_in_67,dangling_wire_437,demux_data_in_66,dangling_wire_438,demux_data_in_65,dangling_wire_439,demux_data_in_64}),
            .RADDR({dangling_wire_440,dangling_wire_441,N__18106,N__16189,N__16405,N__16606,N__14791,N__15019,N__15205,N__15433,N__15646}),
            .WADDR({dangling_wire_442,dangling_wire_443,N__18109,N__16207,N__16423,N__16627,N__14806,N__15010,N__15226,N__15436,N__15673}),
            .MASK({dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459}),
            .WDATA({dangling_wire_460,N__13485,dangling_wire_461,N__13663,dangling_wire_462,N__13826,dangling_wire_463,N__12650,dangling_wire_464,N__12779,dangling_wire_465,N__12894,dangling_wire_466,N__13007,dangling_wire_467,N__13125}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26153),
            .WCLKE(N__13270),
            .WCLK(N__27473),
            .WE(N__26149));
    defparam \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \genblk1_genblk1_9__ram_i.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_468,demux_data_in_79,dangling_wire_469,demux_data_in_78,dangling_wire_470,demux_data_in_77,dangling_wire_471,demux_data_in_76,dangling_wire_472,demux_data_in_75,dangling_wire_473,demux_data_in_74,dangling_wire_474,demux_data_in_73,dangling_wire_475,demux_data_in_72}),
            .RADDR({dangling_wire_476,dangling_wire_477,N__18082,N__16164,N__16380,N__16581,N__14766,N__14995,N__15180,N__15409,N__15622}),
            .WADDR({dangling_wire_478,dangling_wire_479,N__18085,N__16183,N__16399,N__16603,N__14782,N__14986,N__15202,N__15412,N__15649}),
            .MASK({dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495}),
            .WDATA({dangling_wire_496,N__13486,dangling_wire_497,N__13664,dangling_wire_498,N__13831,dangling_wire_499,N__12651,dangling_wire_500,N__12784,dangling_wire_501,N__12908,dangling_wire_502,N__13008,dangling_wire_503,N__13126}),
            .RCLKE(),
            .RCLK(\INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net ),
            .RE(N__26154),
            .WCLKE(N__11173),
            .WCLK(N__27488),
            .WE(N__26195));
    IO_PAD_OD reset_n_input_iopad_od (
            .OE(N__28196),
            .DIN(N__28195),
            .DOUT(N__28194),
            .PACKAGEPIN(reset_n_in));
    defparam reset_n_input_preio.PIN_TYPE=6'b000001;
    defparam reset_n_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO reset_n_input_preio (
            .PADOEN(N__28196),
            .PADOUT(N__28195),
            .PADIN(N__28194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(reset_n),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD_OD clk_spi_input_iopad_od (
            .OE(N__28187),
            .DIN(N__28186),
            .DOUT(N__28185),
            .PACKAGEPIN(clk_spi_in));
    defparam clk_spi_input_preio.PIN_TYPE=6'b000001;
    defparam clk_spi_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO clk_spi_input_preio (
            .PADOEN(N__28187),
            .PADOUT(N__28186),
            .PADIN(N__28185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_spi),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD_OD miso_output_iopad_od (
            .OE(N__28178),
            .DIN(N__28177),
            .DOUT(N__28176),
            .PACKAGEPIN(miso_out));
    defparam miso_output_preio.PIN_TYPE=6'b011001;
    defparam miso_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO miso_output_preio (
            .PADOEN(N__28178),
            .PADOUT(N__28177),
            .PADIN(N__28176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD_OD cs_n_input_iopad_od (
            .OE(N__28169),
            .DIN(N__28168),
            .DOUT(N__28167),
            .PACKAGEPIN(cs_n_in));
    defparam cs_n_input_preio.PIN_TYPE=6'b000001;
    defparam cs_n_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO cs_n_input_preio (
            .PADOEN(N__28169),
            .PADOUT(N__28168),
            .PADIN(N__28167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(cs_n),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD_OD mosi_input_iopad_od (
            .OE(N__28160),
            .DIN(N__28159),
            .DOUT(N__28158),
            .PACKAGEPIN(mosi_in));
    defparam mosi_input_preio.PIN_TYPE=6'b000001;
    defparam mosi_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO mosi_input_preio (
            .PADOEN(N__28160),
            .PADOUT(N__28159),
            .PADIN(N__28158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(mosi),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_output_iopad (
            .OE(N__28151),
            .DIN(N__28150),
            .DOUT(N__28149),
            .PACKAGEPIN(led_out));
    defparam led_output_preio.PIN_TYPE=6'b011000;
    defparam led_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO led_output_preio (
            .PADOEN(N__28151),
            .PADOUT(N__28150),
            .PADIN(N__28149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24811),
            .INPUTCLK(GNDG0),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__6847 (
            .O(N__28132),
            .I(N__28129));
    InMux I__6846 (
            .O(N__28129),
            .I(N__28126));
    LocalMux I__6845 (
            .O(N__28126),
            .I(\ws2812.rgb_counter_0_sqmuxa_0_a2_0_1 ));
    InMux I__6844 (
            .O(N__28123),
            .I(N__28119));
    CascadeMux I__6843 (
            .O(N__28122),
            .I(N__28103));
    LocalMux I__6842 (
            .O(N__28119),
            .I(N__28100));
    InMux I__6841 (
            .O(N__28118),
            .I(N__28097));
    InMux I__6840 (
            .O(N__28117),
            .I(N__28088));
    InMux I__6839 (
            .O(N__28116),
            .I(N__28088));
    InMux I__6838 (
            .O(N__28115),
            .I(N__28088));
    InMux I__6837 (
            .O(N__28114),
            .I(N__28088));
    InMux I__6836 (
            .O(N__28113),
            .I(N__28083));
    InMux I__6835 (
            .O(N__28112),
            .I(N__28083));
    InMux I__6834 (
            .O(N__28111),
            .I(N__28078));
    InMux I__6833 (
            .O(N__28110),
            .I(N__28078));
    InMux I__6832 (
            .O(N__28109),
            .I(N__28073));
    InMux I__6831 (
            .O(N__28108),
            .I(N__28073));
    InMux I__6830 (
            .O(N__28107),
            .I(N__28068));
    InMux I__6829 (
            .O(N__28106),
            .I(N__28068));
    InMux I__6828 (
            .O(N__28103),
            .I(N__28065));
    Odrv4 I__6827 (
            .O(N__28100),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6826 (
            .O(N__28097),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6825 (
            .O(N__28088),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6824 (
            .O(N__28083),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6823 (
            .O(N__28078),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6822 (
            .O(N__28073),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6821 (
            .O(N__28068),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    LocalMux I__6820 (
            .O(N__28065),
            .I(\ws2812.rgb_counterZ0Z_2 ));
    CascadeMux I__6819 (
            .O(N__28048),
            .I(N__28045));
    InMux I__6818 (
            .O(N__28045),
            .I(N__28042));
    LocalMux I__6817 (
            .O(N__28042),
            .I(\ws2812.rgb_counter_RNI2AOD3Z0Z_2 ));
    InMux I__6816 (
            .O(N__28039),
            .I(N__28036));
    LocalMux I__6815 (
            .O(N__28036),
            .I(N__28029));
    InMux I__6814 (
            .O(N__28035),
            .I(N__28026));
    InMux I__6813 (
            .O(N__28034),
            .I(N__28023));
    InMux I__6812 (
            .O(N__28033),
            .I(N__28020));
    InMux I__6811 (
            .O(N__28032),
            .I(N__28017));
    Odrv4 I__6810 (
            .O(N__28029),
            .I(\ws2812.rgb_counterZ0Z_1 ));
    LocalMux I__6809 (
            .O(N__28026),
            .I(\ws2812.rgb_counterZ0Z_1 ));
    LocalMux I__6808 (
            .O(N__28023),
            .I(\ws2812.rgb_counterZ0Z_1 ));
    LocalMux I__6807 (
            .O(N__28020),
            .I(\ws2812.rgb_counterZ0Z_1 ));
    LocalMux I__6806 (
            .O(N__28017),
            .I(\ws2812.rgb_counterZ0Z_1 ));
    CascadeMux I__6805 (
            .O(N__28006),
            .I(N__28003));
    InMux I__6804 (
            .O(N__28003),
            .I(N__28000));
    LocalMux I__6803 (
            .O(N__28000),
            .I(\ws2812.rgb_counter_RNI19OD3Z0Z_1 ));
    InMux I__6802 (
            .O(N__27997),
            .I(N__27991));
    InMux I__6801 (
            .O(N__27996),
            .I(N__27988));
    InMux I__6800 (
            .O(N__27995),
            .I(N__27985));
    InMux I__6799 (
            .O(N__27994),
            .I(N__27982));
    LocalMux I__6798 (
            .O(N__27991),
            .I(N__27979));
    LocalMux I__6797 (
            .O(N__27988),
            .I(N__27976));
    LocalMux I__6796 (
            .O(N__27985),
            .I(N__27973));
    LocalMux I__6795 (
            .O(N__27982),
            .I(N__27970));
    Span4Mux_v I__6794 (
            .O(N__27979),
            .I(N__27967));
    Span4Mux_v I__6793 (
            .O(N__27976),
            .I(N__27964));
    Span4Mux_s3_h I__6792 (
            .O(N__27973),
            .I(N__27961));
    Span4Mux_v I__6791 (
            .O(N__27970),
            .I(N__27958));
    Odrv4 I__6790 (
            .O(N__27967),
            .I(\ws2812.rgb_counterZ0Z_3 ));
    Odrv4 I__6789 (
            .O(N__27964),
            .I(\ws2812.rgb_counterZ0Z_3 ));
    Odrv4 I__6788 (
            .O(N__27961),
            .I(\ws2812.rgb_counterZ0Z_3 ));
    Odrv4 I__6787 (
            .O(N__27958),
            .I(\ws2812.rgb_counterZ0Z_3 ));
    CascadeMux I__6786 (
            .O(N__27949),
            .I(N__27946));
    InMux I__6785 (
            .O(N__27946),
            .I(N__27943));
    LocalMux I__6784 (
            .O(N__27943),
            .I(\ws2812.rgb_counter_RNI3BOD3Z0Z_3 ));
    InMux I__6783 (
            .O(N__27940),
            .I(N__27937));
    LocalMux I__6782 (
            .O(N__27937),
            .I(N__27928));
    InMux I__6781 (
            .O(N__27936),
            .I(N__27925));
    InMux I__6780 (
            .O(N__27935),
            .I(N__27922));
    InMux I__6779 (
            .O(N__27934),
            .I(N__27917));
    InMux I__6778 (
            .O(N__27933),
            .I(N__27917));
    InMux I__6777 (
            .O(N__27932),
            .I(N__27912));
    InMux I__6776 (
            .O(N__27931),
            .I(N__27912));
    Span4Mux_v I__6775 (
            .O(N__27928),
            .I(N__27908));
    LocalMux I__6774 (
            .O(N__27925),
            .I(N__27903));
    LocalMux I__6773 (
            .O(N__27922),
            .I(N__27903));
    LocalMux I__6772 (
            .O(N__27917),
            .I(N__27900));
    LocalMux I__6771 (
            .O(N__27912),
            .I(N__27897));
    InMux I__6770 (
            .O(N__27911),
            .I(N__27894));
    Span4Mux_s0_h I__6769 (
            .O(N__27908),
            .I(N__27889));
    Span4Mux_v I__6768 (
            .O(N__27903),
            .I(N__27889));
    Span4Mux_v I__6767 (
            .O(N__27900),
            .I(N__27886));
    Span4Mux_s3_h I__6766 (
            .O(N__27897),
            .I(N__27883));
    LocalMux I__6765 (
            .O(N__27894),
            .I(\ws2812.rgb_counterZ0Z_0 ));
    Odrv4 I__6764 (
            .O(N__27889),
            .I(\ws2812.rgb_counterZ0Z_0 ));
    Odrv4 I__6763 (
            .O(N__27886),
            .I(\ws2812.rgb_counterZ0Z_0 ));
    Odrv4 I__6762 (
            .O(N__27883),
            .I(\ws2812.rgb_counterZ0Z_0 ));
    CascadeMux I__6761 (
            .O(N__27874),
            .I(N__27871));
    InMux I__6760 (
            .O(N__27871),
            .I(N__27868));
    LocalMux I__6759 (
            .O(N__27868),
            .I(\ws2812.un1_rgb_counter_cry_0_c_RNOZ0 ));
    CascadeMux I__6758 (
            .O(N__27865),
            .I(N__27852));
    InMux I__6757 (
            .O(N__27864),
            .I(N__27845));
    InMux I__6756 (
            .O(N__27863),
            .I(N__27845));
    InMux I__6755 (
            .O(N__27862),
            .I(N__27845));
    InMux I__6754 (
            .O(N__27861),
            .I(N__27842));
    InMux I__6753 (
            .O(N__27860),
            .I(N__27831));
    InMux I__6752 (
            .O(N__27859),
            .I(N__27831));
    InMux I__6751 (
            .O(N__27858),
            .I(N__27831));
    InMux I__6750 (
            .O(N__27857),
            .I(N__27831));
    InMux I__6749 (
            .O(N__27856),
            .I(N__27831));
    InMux I__6748 (
            .O(N__27855),
            .I(N__27825));
    InMux I__6747 (
            .O(N__27852),
            .I(N__27822));
    LocalMux I__6746 (
            .O(N__27845),
            .I(N__27819));
    LocalMux I__6745 (
            .O(N__27842),
            .I(N__27814));
    LocalMux I__6744 (
            .O(N__27831),
            .I(N__27814));
    InMux I__6743 (
            .O(N__27830),
            .I(N__27809));
    InMux I__6742 (
            .O(N__27829),
            .I(N__27809));
    InMux I__6741 (
            .O(N__27828),
            .I(N__27806));
    LocalMux I__6740 (
            .O(N__27825),
            .I(N__27801));
    LocalMux I__6739 (
            .O(N__27822),
            .I(N__27801));
    Span4Mux_v I__6738 (
            .O(N__27819),
            .I(N__27796));
    Span4Mux_v I__6737 (
            .O(N__27814),
            .I(N__27796));
    LocalMux I__6736 (
            .O(N__27809),
            .I(\ws2812.N_106 ));
    LocalMux I__6735 (
            .O(N__27806),
            .I(\ws2812.N_106 ));
    Odrv12 I__6734 (
            .O(N__27801),
            .I(\ws2812.N_106 ));
    Odrv4 I__6733 (
            .O(N__27796),
            .I(\ws2812.N_106 ));
    InMux I__6732 (
            .O(N__27787),
            .I(N__27783));
    InMux I__6731 (
            .O(N__27786),
            .I(N__27780));
    LocalMux I__6730 (
            .O(N__27783),
            .I(N__27777));
    LocalMux I__6729 (
            .O(N__27780),
            .I(N__27774));
    Span4Mux_s0_h I__6728 (
            .O(N__27777),
            .I(N__27771));
    Span12Mux_s7_v I__6727 (
            .O(N__27774),
            .I(N__27766));
    Span4Mux_h I__6726 (
            .O(N__27771),
            .I(N__27763));
    InMux I__6725 (
            .O(N__27770),
            .I(N__27758));
    InMux I__6724 (
            .O(N__27769),
            .I(N__27758));
    Odrv12 I__6723 (
            .O(N__27766),
            .I(send_leds_n));
    Odrv4 I__6722 (
            .O(N__27763),
            .I(send_leds_n));
    LocalMux I__6721 (
            .O(N__27758),
            .I(send_leds_n));
    CascadeMux I__6720 (
            .O(N__27751),
            .I(N__27738));
    InMux I__6719 (
            .O(N__27750),
            .I(N__27727));
    InMux I__6718 (
            .O(N__27749),
            .I(N__27727));
    CascadeMux I__6717 (
            .O(N__27748),
            .I(N__27724));
    CascadeMux I__6716 (
            .O(N__27747),
            .I(N__27720));
    CascadeMux I__6715 (
            .O(N__27746),
            .I(N__27716));
    CascadeMux I__6714 (
            .O(N__27745),
            .I(N__27712));
    CascadeMux I__6713 (
            .O(N__27744),
            .I(N__27708));
    CascadeMux I__6712 (
            .O(N__27743),
            .I(N__27705));
    CascadeMux I__6711 (
            .O(N__27742),
            .I(N__27702));
    InMux I__6710 (
            .O(N__27741),
            .I(N__27697));
    InMux I__6709 (
            .O(N__27738),
            .I(N__27693));
    InMux I__6708 (
            .O(N__27737),
            .I(N__27680));
    InMux I__6707 (
            .O(N__27736),
            .I(N__27680));
    InMux I__6706 (
            .O(N__27735),
            .I(N__27680));
    InMux I__6705 (
            .O(N__27734),
            .I(N__27680));
    InMux I__6704 (
            .O(N__27733),
            .I(N__27680));
    InMux I__6703 (
            .O(N__27732),
            .I(N__27680));
    LocalMux I__6702 (
            .O(N__27727),
            .I(N__27676));
    InMux I__6701 (
            .O(N__27724),
            .I(N__27661));
    InMux I__6700 (
            .O(N__27723),
            .I(N__27661));
    InMux I__6699 (
            .O(N__27720),
            .I(N__27661));
    InMux I__6698 (
            .O(N__27719),
            .I(N__27661));
    InMux I__6697 (
            .O(N__27716),
            .I(N__27661));
    InMux I__6696 (
            .O(N__27715),
            .I(N__27661));
    InMux I__6695 (
            .O(N__27712),
            .I(N__27661));
    InMux I__6694 (
            .O(N__27711),
            .I(N__27658));
    InMux I__6693 (
            .O(N__27708),
            .I(N__27647));
    InMux I__6692 (
            .O(N__27705),
            .I(N__27647));
    InMux I__6691 (
            .O(N__27702),
            .I(N__27647));
    InMux I__6690 (
            .O(N__27701),
            .I(N__27647));
    InMux I__6689 (
            .O(N__27700),
            .I(N__27647));
    LocalMux I__6688 (
            .O(N__27697),
            .I(N__27644));
    InMux I__6687 (
            .O(N__27696),
            .I(N__27641));
    LocalMux I__6686 (
            .O(N__27693),
            .I(N__27636));
    LocalMux I__6685 (
            .O(N__27680),
            .I(N__27636));
    InMux I__6684 (
            .O(N__27679),
            .I(N__27633));
    Span12Mux_s5_v I__6683 (
            .O(N__27676),
            .I(N__27628));
    LocalMux I__6682 (
            .O(N__27661),
            .I(N__27628));
    LocalMux I__6681 (
            .O(N__27658),
            .I(N__27621));
    LocalMux I__6680 (
            .O(N__27647),
            .I(N__27621));
    Span4Mux_h I__6679 (
            .O(N__27644),
            .I(N__27621));
    LocalMux I__6678 (
            .O(N__27641),
            .I(N__27616));
    Span4Mux_h I__6677 (
            .O(N__27636),
            .I(N__27616));
    LocalMux I__6676 (
            .O(N__27633),
            .I(\ws2812.stateZ0Z_0 ));
    Odrv12 I__6675 (
            .O(N__27628),
            .I(\ws2812.stateZ0Z_0 ));
    Odrv4 I__6674 (
            .O(N__27621),
            .I(\ws2812.stateZ0Z_0 ));
    Odrv4 I__6673 (
            .O(N__27616),
            .I(\ws2812.stateZ0Z_0 ));
    CascadeMux I__6672 (
            .O(N__27607),
            .I(N__27604));
    InMux I__6671 (
            .O(N__27604),
            .I(N__27601));
    LocalMux I__6670 (
            .O(N__27601),
            .I(N__27597));
    InMux I__6669 (
            .O(N__27600),
            .I(N__27594));
    Span4Mux_v I__6668 (
            .O(N__27597),
            .I(N__27589));
    LocalMux I__6667 (
            .O(N__27594),
            .I(N__27589));
    Span4Mux_h I__6666 (
            .O(N__27589),
            .I(N__27585));
    InMux I__6665 (
            .O(N__27588),
            .I(N__27582));
    Odrv4 I__6664 (
            .O(N__27585),
            .I(\ws2812.N_228 ));
    LocalMux I__6663 (
            .O(N__27582),
            .I(\ws2812.N_228 ));
    InMux I__6662 (
            .O(N__27577),
            .I(N__27569));
    InMux I__6661 (
            .O(N__27576),
            .I(N__27569));
    InMux I__6660 (
            .O(N__27575),
            .I(N__27566));
    InMux I__6659 (
            .O(N__27574),
            .I(N__27563));
    LocalMux I__6658 (
            .O(N__27569),
            .I(N__27559));
    LocalMux I__6657 (
            .O(N__27566),
            .I(N__27556));
    LocalMux I__6656 (
            .O(N__27563),
            .I(N__27553));
    InMux I__6655 (
            .O(N__27562),
            .I(N__27550));
    Span4Mux_v I__6654 (
            .O(N__27559),
            .I(N__27545));
    Span4Mux_h I__6653 (
            .O(N__27556),
            .I(N__27545));
    Span4Mux_h I__6652 (
            .O(N__27553),
            .I(N__27540));
    LocalMux I__6651 (
            .O(N__27550),
            .I(N__27540));
    Odrv4 I__6650 (
            .O(N__27545),
            .I(\ws2812.state_RNIELS35Z0Z_0 ));
    Odrv4 I__6649 (
            .O(N__27540),
            .I(\ws2812.state_RNIELS35Z0Z_0 ));
    InMux I__6648 (
            .O(N__27535),
            .I(N__27532));
    LocalMux I__6647 (
            .O(N__27532),
            .I(N__27529));
    Odrv12 I__6646 (
            .O(N__27529),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_6 ));
    InMux I__6645 (
            .O(N__27526),
            .I(N__27523));
    LocalMux I__6644 (
            .O(N__27523),
            .I(rgb_data_out_6));
    ClkMux I__6643 (
            .O(N__27520),
            .I(N__27214));
    ClkMux I__6642 (
            .O(N__27519),
            .I(N__27214));
    ClkMux I__6641 (
            .O(N__27518),
            .I(N__27214));
    ClkMux I__6640 (
            .O(N__27517),
            .I(N__27214));
    ClkMux I__6639 (
            .O(N__27516),
            .I(N__27214));
    ClkMux I__6638 (
            .O(N__27515),
            .I(N__27214));
    ClkMux I__6637 (
            .O(N__27514),
            .I(N__27214));
    ClkMux I__6636 (
            .O(N__27513),
            .I(N__27214));
    ClkMux I__6635 (
            .O(N__27512),
            .I(N__27214));
    ClkMux I__6634 (
            .O(N__27511),
            .I(N__27214));
    ClkMux I__6633 (
            .O(N__27510),
            .I(N__27214));
    ClkMux I__6632 (
            .O(N__27509),
            .I(N__27214));
    ClkMux I__6631 (
            .O(N__27508),
            .I(N__27214));
    ClkMux I__6630 (
            .O(N__27507),
            .I(N__27214));
    ClkMux I__6629 (
            .O(N__27506),
            .I(N__27214));
    ClkMux I__6628 (
            .O(N__27505),
            .I(N__27214));
    ClkMux I__6627 (
            .O(N__27504),
            .I(N__27214));
    ClkMux I__6626 (
            .O(N__27503),
            .I(N__27214));
    ClkMux I__6625 (
            .O(N__27502),
            .I(N__27214));
    ClkMux I__6624 (
            .O(N__27501),
            .I(N__27214));
    ClkMux I__6623 (
            .O(N__27500),
            .I(N__27214));
    ClkMux I__6622 (
            .O(N__27499),
            .I(N__27214));
    ClkMux I__6621 (
            .O(N__27498),
            .I(N__27214));
    ClkMux I__6620 (
            .O(N__27497),
            .I(N__27214));
    ClkMux I__6619 (
            .O(N__27496),
            .I(N__27214));
    ClkMux I__6618 (
            .O(N__27495),
            .I(N__27214));
    ClkMux I__6617 (
            .O(N__27494),
            .I(N__27214));
    ClkMux I__6616 (
            .O(N__27493),
            .I(N__27214));
    ClkMux I__6615 (
            .O(N__27492),
            .I(N__27214));
    ClkMux I__6614 (
            .O(N__27491),
            .I(N__27214));
    ClkMux I__6613 (
            .O(N__27490),
            .I(N__27214));
    ClkMux I__6612 (
            .O(N__27489),
            .I(N__27214));
    ClkMux I__6611 (
            .O(N__27488),
            .I(N__27214));
    ClkMux I__6610 (
            .O(N__27487),
            .I(N__27214));
    ClkMux I__6609 (
            .O(N__27486),
            .I(N__27214));
    ClkMux I__6608 (
            .O(N__27485),
            .I(N__27214));
    ClkMux I__6607 (
            .O(N__27484),
            .I(N__27214));
    ClkMux I__6606 (
            .O(N__27483),
            .I(N__27214));
    ClkMux I__6605 (
            .O(N__27482),
            .I(N__27214));
    ClkMux I__6604 (
            .O(N__27481),
            .I(N__27214));
    ClkMux I__6603 (
            .O(N__27480),
            .I(N__27214));
    ClkMux I__6602 (
            .O(N__27479),
            .I(N__27214));
    ClkMux I__6601 (
            .O(N__27478),
            .I(N__27214));
    ClkMux I__6600 (
            .O(N__27477),
            .I(N__27214));
    ClkMux I__6599 (
            .O(N__27476),
            .I(N__27214));
    ClkMux I__6598 (
            .O(N__27475),
            .I(N__27214));
    ClkMux I__6597 (
            .O(N__27474),
            .I(N__27214));
    ClkMux I__6596 (
            .O(N__27473),
            .I(N__27214));
    ClkMux I__6595 (
            .O(N__27472),
            .I(N__27214));
    ClkMux I__6594 (
            .O(N__27471),
            .I(N__27214));
    ClkMux I__6593 (
            .O(N__27470),
            .I(N__27214));
    ClkMux I__6592 (
            .O(N__27469),
            .I(N__27214));
    ClkMux I__6591 (
            .O(N__27468),
            .I(N__27214));
    ClkMux I__6590 (
            .O(N__27467),
            .I(N__27214));
    ClkMux I__6589 (
            .O(N__27466),
            .I(N__27214));
    ClkMux I__6588 (
            .O(N__27465),
            .I(N__27214));
    ClkMux I__6587 (
            .O(N__27464),
            .I(N__27214));
    ClkMux I__6586 (
            .O(N__27463),
            .I(N__27214));
    ClkMux I__6585 (
            .O(N__27462),
            .I(N__27214));
    ClkMux I__6584 (
            .O(N__27461),
            .I(N__27214));
    ClkMux I__6583 (
            .O(N__27460),
            .I(N__27214));
    ClkMux I__6582 (
            .O(N__27459),
            .I(N__27214));
    ClkMux I__6581 (
            .O(N__27458),
            .I(N__27214));
    ClkMux I__6580 (
            .O(N__27457),
            .I(N__27214));
    ClkMux I__6579 (
            .O(N__27456),
            .I(N__27214));
    ClkMux I__6578 (
            .O(N__27455),
            .I(N__27214));
    ClkMux I__6577 (
            .O(N__27454),
            .I(N__27214));
    ClkMux I__6576 (
            .O(N__27453),
            .I(N__27214));
    ClkMux I__6575 (
            .O(N__27452),
            .I(N__27214));
    ClkMux I__6574 (
            .O(N__27451),
            .I(N__27214));
    ClkMux I__6573 (
            .O(N__27450),
            .I(N__27214));
    ClkMux I__6572 (
            .O(N__27449),
            .I(N__27214));
    ClkMux I__6571 (
            .O(N__27448),
            .I(N__27214));
    ClkMux I__6570 (
            .O(N__27447),
            .I(N__27214));
    ClkMux I__6569 (
            .O(N__27446),
            .I(N__27214));
    ClkMux I__6568 (
            .O(N__27445),
            .I(N__27214));
    ClkMux I__6567 (
            .O(N__27444),
            .I(N__27214));
    ClkMux I__6566 (
            .O(N__27443),
            .I(N__27214));
    ClkMux I__6565 (
            .O(N__27442),
            .I(N__27214));
    ClkMux I__6564 (
            .O(N__27441),
            .I(N__27214));
    ClkMux I__6563 (
            .O(N__27440),
            .I(N__27214));
    ClkMux I__6562 (
            .O(N__27439),
            .I(N__27214));
    ClkMux I__6561 (
            .O(N__27438),
            .I(N__27214));
    ClkMux I__6560 (
            .O(N__27437),
            .I(N__27214));
    ClkMux I__6559 (
            .O(N__27436),
            .I(N__27214));
    ClkMux I__6558 (
            .O(N__27435),
            .I(N__27214));
    ClkMux I__6557 (
            .O(N__27434),
            .I(N__27214));
    ClkMux I__6556 (
            .O(N__27433),
            .I(N__27214));
    ClkMux I__6555 (
            .O(N__27432),
            .I(N__27214));
    ClkMux I__6554 (
            .O(N__27431),
            .I(N__27214));
    ClkMux I__6553 (
            .O(N__27430),
            .I(N__27214));
    ClkMux I__6552 (
            .O(N__27429),
            .I(N__27214));
    ClkMux I__6551 (
            .O(N__27428),
            .I(N__27214));
    ClkMux I__6550 (
            .O(N__27427),
            .I(N__27214));
    ClkMux I__6549 (
            .O(N__27426),
            .I(N__27214));
    ClkMux I__6548 (
            .O(N__27425),
            .I(N__27214));
    ClkMux I__6547 (
            .O(N__27424),
            .I(N__27214));
    ClkMux I__6546 (
            .O(N__27423),
            .I(N__27214));
    ClkMux I__6545 (
            .O(N__27422),
            .I(N__27214));
    ClkMux I__6544 (
            .O(N__27421),
            .I(N__27214));
    ClkMux I__6543 (
            .O(N__27420),
            .I(N__27214));
    ClkMux I__6542 (
            .O(N__27419),
            .I(N__27214));
    GlobalMux I__6541 (
            .O(N__27214),
            .I(N__27211));
    DummyBuf I__6540 (
            .O(N__27211),
            .I(clk_sb));
    InMux I__6539 (
            .O(N__27208),
            .I(N__27201));
    InMux I__6538 (
            .O(N__27207),
            .I(N__27201));
    InMux I__6537 (
            .O(N__27206),
            .I(N__27198));
    LocalMux I__6536 (
            .O(N__27201),
            .I(N__27188));
    LocalMux I__6535 (
            .O(N__27198),
            .I(N__27185));
    CEMux I__6534 (
            .O(N__27197),
            .I(N__27166));
    CEMux I__6533 (
            .O(N__27196),
            .I(N__27166));
    CEMux I__6532 (
            .O(N__27195),
            .I(N__27166));
    CEMux I__6531 (
            .O(N__27194),
            .I(N__27166));
    CEMux I__6530 (
            .O(N__27193),
            .I(N__27166));
    CEMux I__6529 (
            .O(N__27192),
            .I(N__27166));
    CEMux I__6528 (
            .O(N__27191),
            .I(N__27166));
    Glb2LocalMux I__6527 (
            .O(N__27188),
            .I(N__27166));
    Glb2LocalMux I__6526 (
            .O(N__27185),
            .I(N__27166));
    GlobalMux I__6525 (
            .O(N__27166),
            .I(N__27163));
    gio2CtrlBuf I__6524 (
            .O(N__27163),
            .I(\sb_translator_1.state_leds_2_sqmuxa_g ));
    CascadeMux I__6523 (
            .O(N__27160),
            .I(N__27154));
    InMux I__6522 (
            .O(N__27159),
            .I(N__27150));
    InMux I__6521 (
            .O(N__27158),
            .I(N__27143));
    InMux I__6520 (
            .O(N__27157),
            .I(N__27143));
    InMux I__6519 (
            .O(N__27154),
            .I(N__27143));
    InMux I__6518 (
            .O(N__27153),
            .I(N__27140));
    LocalMux I__6517 (
            .O(N__27150),
            .I(N__27120));
    LocalMux I__6516 (
            .O(N__27143),
            .I(N__27117));
    LocalMux I__6515 (
            .O(N__27140),
            .I(N__27104));
    SRMux I__6514 (
            .O(N__27139),
            .I(N__26920));
    SRMux I__6513 (
            .O(N__27138),
            .I(N__26920));
    SRMux I__6512 (
            .O(N__27137),
            .I(N__26920));
    SRMux I__6511 (
            .O(N__27136),
            .I(N__26920));
    SRMux I__6510 (
            .O(N__27135),
            .I(N__26920));
    SRMux I__6509 (
            .O(N__27134),
            .I(N__26920));
    SRMux I__6508 (
            .O(N__27133),
            .I(N__26920));
    SRMux I__6507 (
            .O(N__27132),
            .I(N__26920));
    SRMux I__6506 (
            .O(N__27131),
            .I(N__26920));
    SRMux I__6505 (
            .O(N__27130),
            .I(N__26920));
    SRMux I__6504 (
            .O(N__27129),
            .I(N__26920));
    SRMux I__6503 (
            .O(N__27128),
            .I(N__26920));
    SRMux I__6502 (
            .O(N__27127),
            .I(N__26920));
    SRMux I__6501 (
            .O(N__27126),
            .I(N__26920));
    SRMux I__6500 (
            .O(N__27125),
            .I(N__26920));
    SRMux I__6499 (
            .O(N__27124),
            .I(N__26920));
    SRMux I__6498 (
            .O(N__27123),
            .I(N__26920));
    Glb2LocalMux I__6497 (
            .O(N__27120),
            .I(N__26920));
    Glb2LocalMux I__6496 (
            .O(N__27117),
            .I(N__26920));
    SRMux I__6495 (
            .O(N__27116),
            .I(N__26920));
    SRMux I__6494 (
            .O(N__27115),
            .I(N__26920));
    SRMux I__6493 (
            .O(N__27114),
            .I(N__26920));
    SRMux I__6492 (
            .O(N__27113),
            .I(N__26920));
    SRMux I__6491 (
            .O(N__27112),
            .I(N__26920));
    SRMux I__6490 (
            .O(N__27111),
            .I(N__26920));
    SRMux I__6489 (
            .O(N__27110),
            .I(N__26920));
    SRMux I__6488 (
            .O(N__27109),
            .I(N__26920));
    SRMux I__6487 (
            .O(N__27108),
            .I(N__26920));
    SRMux I__6486 (
            .O(N__27107),
            .I(N__26920));
    Glb2LocalMux I__6485 (
            .O(N__27104),
            .I(N__26920));
    SRMux I__6484 (
            .O(N__27103),
            .I(N__26920));
    SRMux I__6483 (
            .O(N__27102),
            .I(N__26920));
    SRMux I__6482 (
            .O(N__27101),
            .I(N__26920));
    SRMux I__6481 (
            .O(N__27100),
            .I(N__26920));
    SRMux I__6480 (
            .O(N__27099),
            .I(N__26920));
    SRMux I__6479 (
            .O(N__27098),
            .I(N__26920));
    SRMux I__6478 (
            .O(N__27097),
            .I(N__26920));
    SRMux I__6477 (
            .O(N__27096),
            .I(N__26920));
    SRMux I__6476 (
            .O(N__27095),
            .I(N__26920));
    SRMux I__6475 (
            .O(N__27094),
            .I(N__26920));
    SRMux I__6474 (
            .O(N__27093),
            .I(N__26920));
    SRMux I__6473 (
            .O(N__27092),
            .I(N__26920));
    SRMux I__6472 (
            .O(N__27091),
            .I(N__26920));
    SRMux I__6471 (
            .O(N__27090),
            .I(N__26920));
    SRMux I__6470 (
            .O(N__27089),
            .I(N__26920));
    SRMux I__6469 (
            .O(N__27088),
            .I(N__26920));
    SRMux I__6468 (
            .O(N__27087),
            .I(N__26920));
    SRMux I__6467 (
            .O(N__27086),
            .I(N__26920));
    SRMux I__6466 (
            .O(N__27085),
            .I(N__26920));
    SRMux I__6465 (
            .O(N__27084),
            .I(N__26920));
    SRMux I__6464 (
            .O(N__27083),
            .I(N__26920));
    SRMux I__6463 (
            .O(N__27082),
            .I(N__26920));
    SRMux I__6462 (
            .O(N__27081),
            .I(N__26920));
    SRMux I__6461 (
            .O(N__27080),
            .I(N__26920));
    SRMux I__6460 (
            .O(N__27079),
            .I(N__26920));
    SRMux I__6459 (
            .O(N__27078),
            .I(N__26920));
    SRMux I__6458 (
            .O(N__27077),
            .I(N__26920));
    SRMux I__6457 (
            .O(N__27076),
            .I(N__26920));
    SRMux I__6456 (
            .O(N__27075),
            .I(N__26920));
    SRMux I__6455 (
            .O(N__27074),
            .I(N__26920));
    SRMux I__6454 (
            .O(N__27073),
            .I(N__26920));
    SRMux I__6453 (
            .O(N__27072),
            .I(N__26920));
    SRMux I__6452 (
            .O(N__27071),
            .I(N__26920));
    SRMux I__6451 (
            .O(N__27070),
            .I(N__26920));
    SRMux I__6450 (
            .O(N__27069),
            .I(N__26920));
    SRMux I__6449 (
            .O(N__27068),
            .I(N__26920));
    SRMux I__6448 (
            .O(N__27067),
            .I(N__26920));
    SRMux I__6447 (
            .O(N__27066),
            .I(N__26920));
    SRMux I__6446 (
            .O(N__27065),
            .I(N__26920));
    SRMux I__6445 (
            .O(N__27064),
            .I(N__26920));
    SRMux I__6444 (
            .O(N__27063),
            .I(N__26920));
    GlobalMux I__6443 (
            .O(N__26920),
            .I(N__26917));
    gio2CtrlBuf I__6442 (
            .O(N__26917),
            .I(reset_n_i_g));
    InMux I__6441 (
            .O(N__26914),
            .I(N__26911));
    LocalMux I__6440 (
            .O(N__26911),
            .I(N__26908));
    Odrv4 I__6439 (
            .O(N__26908),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_22 ));
    InMux I__6438 (
            .O(N__26905),
            .I(N__26901));
    InMux I__6437 (
            .O(N__26904),
            .I(N__26891));
    LocalMux I__6436 (
            .O(N__26901),
            .I(N__26888));
    InMux I__6435 (
            .O(N__26900),
            .I(N__26873));
    InMux I__6434 (
            .O(N__26899),
            .I(N__26873));
    InMux I__6433 (
            .O(N__26898),
            .I(N__26873));
    InMux I__6432 (
            .O(N__26897),
            .I(N__26873));
    InMux I__6431 (
            .O(N__26896),
            .I(N__26873));
    InMux I__6430 (
            .O(N__26895),
            .I(N__26873));
    InMux I__6429 (
            .O(N__26894),
            .I(N__26873));
    LocalMux I__6428 (
            .O(N__26891),
            .I(N__26869));
    Span4Mux_v I__6427 (
            .O(N__26888),
            .I(N__26864));
    LocalMux I__6426 (
            .O(N__26873),
            .I(N__26864));
    InMux I__6425 (
            .O(N__26872),
            .I(N__26855));
    Span4Mux_s2_h I__6424 (
            .O(N__26869),
            .I(N__26850));
    Span4Mux_h I__6423 (
            .O(N__26864),
            .I(N__26850));
    InMux I__6422 (
            .O(N__26863),
            .I(N__26837));
    InMux I__6421 (
            .O(N__26862),
            .I(N__26837));
    InMux I__6420 (
            .O(N__26861),
            .I(N__26837));
    InMux I__6419 (
            .O(N__26860),
            .I(N__26837));
    InMux I__6418 (
            .O(N__26859),
            .I(N__26837));
    InMux I__6417 (
            .O(N__26858),
            .I(N__26837));
    LocalMux I__6416 (
            .O(N__26855),
            .I(\ws2812.N_105 ));
    Odrv4 I__6415 (
            .O(N__26850),
            .I(\ws2812.N_105 ));
    LocalMux I__6414 (
            .O(N__26837),
            .I(\ws2812.N_105 ));
    InMux I__6413 (
            .O(N__26830),
            .I(N__26827));
    LocalMux I__6412 (
            .O(N__26827),
            .I(N__26824));
    Odrv4 I__6411 (
            .O(N__26824),
            .I(rgb_data_out_23));
    CascadeMux I__6410 (
            .O(N__26821),
            .I(\ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_ ));
    InMux I__6409 (
            .O(N__26818),
            .I(N__26815));
    LocalMux I__6408 (
            .O(N__26815),
            .I(\ws2812.N_117 ));
    InMux I__6407 (
            .O(N__26812),
            .I(N__26809));
    LocalMux I__6406 (
            .O(N__26809),
            .I(N__26806));
    Span4Mux_v I__6405 (
            .O(N__26806),
            .I(N__26803));
    Odrv4 I__6404 (
            .O(N__26803),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_3 ));
    InMux I__6403 (
            .O(N__26800),
            .I(N__26797));
    LocalMux I__6402 (
            .O(N__26797),
            .I(rgb_data_out_3));
    InMux I__6401 (
            .O(N__26794),
            .I(N__26791));
    LocalMux I__6400 (
            .O(N__26791),
            .I(N__26788));
    Span4Mux_v I__6399 (
            .O(N__26788),
            .I(N__26785));
    Odrv4 I__6398 (
            .O(N__26785),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_19 ));
    CascadeMux I__6397 (
            .O(N__26782),
            .I(N__26779));
    InMux I__6396 (
            .O(N__26779),
            .I(N__26776));
    LocalMux I__6395 (
            .O(N__26776),
            .I(rgb_data_out_19));
    InMux I__6394 (
            .O(N__26773),
            .I(N__26770));
    LocalMux I__6393 (
            .O(N__26770),
            .I(N__26767));
    Span12Mux_s4_h I__6392 (
            .O(N__26767),
            .I(N__26764));
    Odrv12 I__6391 (
            .O(N__26764),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_7 ));
    InMux I__6390 (
            .O(N__26761),
            .I(N__26758));
    LocalMux I__6389 (
            .O(N__26758),
            .I(rgb_data_out_7));
    CascadeMux I__6388 (
            .O(N__26755),
            .I(N__26751));
    InMux I__6387 (
            .O(N__26754),
            .I(N__26746));
    InMux I__6386 (
            .O(N__26751),
            .I(N__26741));
    InMux I__6385 (
            .O(N__26750),
            .I(N__26736));
    InMux I__6384 (
            .O(N__26749),
            .I(N__26736));
    LocalMux I__6383 (
            .O(N__26746),
            .I(N__26733));
    InMux I__6382 (
            .O(N__26745),
            .I(N__26728));
    InMux I__6381 (
            .O(N__26744),
            .I(N__26728));
    LocalMux I__6380 (
            .O(N__26741),
            .I(\ws2812.rgb_counter_4 ));
    LocalMux I__6379 (
            .O(N__26736),
            .I(\ws2812.rgb_counter_4 ));
    Odrv4 I__6378 (
            .O(N__26733),
            .I(\ws2812.rgb_counter_4 ));
    LocalMux I__6377 (
            .O(N__26728),
            .I(\ws2812.rgb_counter_4 ));
    CascadeMux I__6376 (
            .O(N__26719),
            .I(N__26716));
    InMux I__6375 (
            .O(N__26716),
            .I(N__26713));
    LocalMux I__6374 (
            .O(N__26713),
            .I(N__26710));
    Odrv4 I__6373 (
            .O(N__26710),
            .I(rgb_data_out_22));
    InMux I__6372 (
            .O(N__26707),
            .I(N__26704));
    LocalMux I__6371 (
            .O(N__26704),
            .I(\ws2812.rgb_data_pmux_6_i_m2_ns_1 ));
    CascadeMux I__6370 (
            .O(N__26701),
            .I(N__26698));
    InMux I__6369 (
            .O(N__26698),
            .I(N__26695));
    LocalMux I__6368 (
            .O(N__26695),
            .I(\ws2812.N_124 ));
    InMux I__6367 (
            .O(N__26692),
            .I(\ws2812.un1_rgb_counter_cry_3 ));
    InMux I__6366 (
            .O(N__26689),
            .I(N__26686));
    LocalMux I__6365 (
            .O(N__26686),
            .I(rgb_data_out_1));
    InMux I__6364 (
            .O(N__26683),
            .I(N__26680));
    LocalMux I__6363 (
            .O(N__26680),
            .I(rgb_data_out_21));
    CascadeMux I__6362 (
            .O(N__26677),
            .I(\ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_ ));
    InMux I__6361 (
            .O(N__26674),
            .I(N__26671));
    LocalMux I__6360 (
            .O(N__26671),
            .I(rgb_data_out_5));
    InMux I__6359 (
            .O(N__26668),
            .I(N__26665));
    LocalMux I__6358 (
            .O(N__26665),
            .I(N__26662));
    Odrv4 I__6357 (
            .O(N__26662),
            .I(\ws2812.N_120 ));
    InMux I__6356 (
            .O(N__26659),
            .I(N__26656));
    LocalMux I__6355 (
            .O(N__26656),
            .I(N__26653));
    Span4Mux_s3_h I__6354 (
            .O(N__26653),
            .I(N__26650));
    Odrv4 I__6353 (
            .O(N__26650),
            .I(rgb_data_out_18));
    InMux I__6352 (
            .O(N__26647),
            .I(N__26644));
    LocalMux I__6351 (
            .O(N__26644),
            .I(N__26641));
    Span4Mux_s2_h I__6350 (
            .O(N__26641),
            .I(N__26638));
    Span4Mux_h I__6349 (
            .O(N__26638),
            .I(N__26635));
    Odrv4 I__6348 (
            .O(N__26635),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_2 ));
    InMux I__6347 (
            .O(N__26632),
            .I(N__26629));
    LocalMux I__6346 (
            .O(N__26629),
            .I(rgb_data_out_2));
    InMux I__6345 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__6344 (
            .O(N__26623),
            .I(N__26620));
    Odrv4 I__6343 (
            .O(N__26620),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_17 ));
    CascadeMux I__6342 (
            .O(N__26617),
            .I(N__26614));
    InMux I__6341 (
            .O(N__26614),
            .I(N__26611));
    LocalMux I__6340 (
            .O(N__26611),
            .I(rgb_data_out_17));
    InMux I__6339 (
            .O(N__26608),
            .I(N__26605));
    LocalMux I__6338 (
            .O(N__26605),
            .I(N__26602));
    Odrv4 I__6337 (
            .O(N__26602),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_23 ));
    InMux I__6336 (
            .O(N__26599),
            .I(N__26596));
    LocalMux I__6335 (
            .O(N__26596),
            .I(N__26593));
    Span4Mux_v I__6334 (
            .O(N__26593),
            .I(N__26590));
    Odrv4 I__6333 (
            .O(N__26590),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_14 ));
    InMux I__6332 (
            .O(N__26587),
            .I(N__26584));
    LocalMux I__6331 (
            .O(N__26584),
            .I(N__26581));
    Odrv4 I__6330 (
            .O(N__26581),
            .I(rgb_data_out_14));
    InMux I__6329 (
            .O(N__26578),
            .I(N__26575));
    LocalMux I__6328 (
            .O(N__26575),
            .I(N__26572));
    Odrv4 I__6327 (
            .O(N__26572),
            .I(\ws2812.data_RNOZ0Z_10 ));
    InMux I__6326 (
            .O(N__26569),
            .I(N__26566));
    LocalMux I__6325 (
            .O(N__26566),
            .I(N__26563));
    Odrv4 I__6324 (
            .O(N__26563),
            .I(\ws2812.data_RNOZ0Z_9 ));
    CascadeMux I__6323 (
            .O(N__26560),
            .I(N__26557));
    InMux I__6322 (
            .O(N__26557),
            .I(N__26554));
    LocalMux I__6321 (
            .O(N__26554),
            .I(N__26551));
    Odrv12 I__6320 (
            .O(N__26551),
            .I(\ws2812.data_RNOZ0Z_8 ));
    InMux I__6319 (
            .O(N__26548),
            .I(N__26545));
    LocalMux I__6318 (
            .O(N__26545),
            .I(\ws2812.N_135 ));
    InMux I__6317 (
            .O(N__26542),
            .I(N__26539));
    LocalMux I__6316 (
            .O(N__26539),
            .I(\ws2812.data_RNOZ0Z_2 ));
    CascadeMux I__6315 (
            .O(N__26536),
            .I(\ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_ ));
    InMux I__6314 (
            .O(N__26533),
            .I(N__26530));
    LocalMux I__6313 (
            .O(N__26530),
            .I(\ws2812.N_115 ));
    CascadeMux I__6312 (
            .O(N__26527),
            .I(N__26524));
    InMux I__6311 (
            .O(N__26524),
            .I(N__26521));
    LocalMux I__6310 (
            .O(N__26521),
            .I(N__26518));
    Odrv12 I__6309 (
            .O(N__26518),
            .I(rgb_data_out_16));
    InMux I__6308 (
            .O(N__26515),
            .I(N__26512));
    LocalMux I__6307 (
            .O(N__26512),
            .I(N__26509));
    Odrv4 I__6306 (
            .O(N__26509),
            .I(rgb_data_out_0));
    InMux I__6305 (
            .O(N__26506),
            .I(N__26503));
    LocalMux I__6304 (
            .O(N__26503),
            .I(N__26500));
    Odrv4 I__6303 (
            .O(N__26500),
            .I(rgb_data_out_20));
    CascadeMux I__6302 (
            .O(N__26497),
            .I(\ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_ ));
    InMux I__6301 (
            .O(N__26494),
            .I(N__26491));
    LocalMux I__6300 (
            .O(N__26491),
            .I(N__26488));
    Odrv4 I__6299 (
            .O(N__26488),
            .I(rgb_data_out_4));
    InMux I__6298 (
            .O(N__26485),
            .I(N__26482));
    LocalMux I__6297 (
            .O(N__26482),
            .I(\ws2812.N_127 ));
    InMux I__6296 (
            .O(N__26479),
            .I(\ws2812.un1_rgb_counter_cry_0 ));
    InMux I__6295 (
            .O(N__26476),
            .I(\ws2812.un1_rgb_counter_cry_1 ));
    InMux I__6294 (
            .O(N__26473),
            .I(N__26470));
    LocalMux I__6293 (
            .O(N__26470),
            .I(N__26467));
    Span4Mux_h I__6292 (
            .O(N__26467),
            .I(N__26464));
    Odrv4 I__6291 (
            .O(N__26464),
            .I(\ws2812.rgb_counter_RNO_0Z0Z_3 ));
    InMux I__6290 (
            .O(N__26461),
            .I(\ws2812.un1_rgb_counter_cry_2 ));
    InMux I__6289 (
            .O(N__26458),
            .I(N__26455));
    LocalMux I__6288 (
            .O(N__26455),
            .I(\ws2812.un6_data_axb_8 ));
    InMux I__6287 (
            .O(N__26452),
            .I(bfn_12_6_0_));
    InMux I__6286 (
            .O(N__26449),
            .I(\ws2812.un6_data_cry_8 ));
    InMux I__6285 (
            .O(N__26446),
            .I(\ws2812.un6_data_cry_9 ));
    InMux I__6284 (
            .O(N__26443),
            .I(N__26440));
    LocalMux I__6283 (
            .O(N__26440),
            .I(N__26437));
    Odrv4 I__6282 (
            .O(N__26437),
            .I(\ws2812.un6_data_axb_11 ));
    InMux I__6281 (
            .O(N__26434),
            .I(\ws2812.un6_data_cry_10 ));
    InMux I__6280 (
            .O(N__26431),
            .I(N__26428));
    LocalMux I__6279 (
            .O(N__26428),
            .I(\ws2812.data_RNOZ0Z_11 ));
    InMux I__6278 (
            .O(N__26425),
            .I(N__26422));
    LocalMux I__6277 (
            .O(N__26422),
            .I(\ws2812.data_RNOZ0Z_12 ));
    CascadeMux I__6276 (
            .O(N__26419),
            .I(N__26416));
    InMux I__6275 (
            .O(N__26416),
            .I(N__26413));
    LocalMux I__6274 (
            .O(N__26413),
            .I(\ws2812.data_RNOZ0Z_13 ));
    InMux I__6273 (
            .O(N__26410),
            .I(\ws2812.un6_data_cry_11 ));
    InMux I__6272 (
            .O(N__26407),
            .I(N__26404));
    LocalMux I__6271 (
            .O(N__26404),
            .I(N__26399));
    InMux I__6270 (
            .O(N__26403),
            .I(N__26396));
    InMux I__6269 (
            .O(N__26402),
            .I(N__26393));
    Span4Mux_v I__6268 (
            .O(N__26399),
            .I(N__26389));
    LocalMux I__6267 (
            .O(N__26396),
            .I(N__26384));
    LocalMux I__6266 (
            .O(N__26393),
            .I(N__26384));
    InMux I__6265 (
            .O(N__26392),
            .I(N__26381));
    Odrv4 I__6264 (
            .O(N__26389),
            .I(\ws2812.bit_counter_10 ));
    Odrv4 I__6263 (
            .O(N__26384),
            .I(\ws2812.bit_counter_10 ));
    LocalMux I__6262 (
            .O(N__26381),
            .I(\ws2812.bit_counter_10 ));
    InMux I__6261 (
            .O(N__26374),
            .I(N__26371));
    LocalMux I__6260 (
            .O(N__26371),
            .I(\ws2812.un6_data_axb_10 ));
    CascadeMux I__6259 (
            .O(N__26368),
            .I(N__26365));
    InMux I__6258 (
            .O(N__26365),
            .I(N__26361));
    CascadeMux I__6257 (
            .O(N__26364),
            .I(N__26358));
    LocalMux I__6256 (
            .O(N__26361),
            .I(N__26355));
    InMux I__6255 (
            .O(N__26358),
            .I(N__26350));
    Span4Mux_h I__6254 (
            .O(N__26355),
            .I(N__26347));
    InMux I__6253 (
            .O(N__26354),
            .I(N__26344));
    InMux I__6252 (
            .O(N__26353),
            .I(N__26341));
    LocalMux I__6251 (
            .O(N__26350),
            .I(N__26338));
    Odrv4 I__6250 (
            .O(N__26347),
            .I(\ws2812.bit_counter_9 ));
    LocalMux I__6249 (
            .O(N__26344),
            .I(\ws2812.bit_counter_9 ));
    LocalMux I__6248 (
            .O(N__26341),
            .I(\ws2812.bit_counter_9 ));
    Odrv4 I__6247 (
            .O(N__26338),
            .I(\ws2812.bit_counter_9 ));
    InMux I__6246 (
            .O(N__26329),
            .I(N__26326));
    LocalMux I__6245 (
            .O(N__26326),
            .I(\ws2812.un6_data_axb_9 ));
    InMux I__6244 (
            .O(N__26323),
            .I(N__26320));
    LocalMux I__6243 (
            .O(N__26320),
            .I(\ws2812.data_RNOZ0Z_6 ));
    InMux I__6242 (
            .O(N__26317),
            .I(N__26314));
    LocalMux I__6241 (
            .O(N__26314),
            .I(\ws2812.data_RNOZ0Z_5 ));
    CascadeMux I__6240 (
            .O(N__26311),
            .I(N__26308));
    InMux I__6239 (
            .O(N__26308),
            .I(N__26305));
    LocalMux I__6238 (
            .O(N__26305),
            .I(\ws2812.data_5_iv_0_47_a2_0_a2_0 ));
    InMux I__6237 (
            .O(N__26302),
            .I(N__26299));
    LocalMux I__6236 (
            .O(N__26299),
            .I(\ws2812.data_5_iv_0_47_a2_0_a2_6_1 ));
    InMux I__6235 (
            .O(N__26296),
            .I(N__26293));
    LocalMux I__6234 (
            .O(N__26293),
            .I(\ws2812.data_5_iv_0_47_a2_0_a2_6 ));
    InMux I__6233 (
            .O(N__26290),
            .I(N__26286));
    InMux I__6232 (
            .O(N__26289),
            .I(N__26283));
    LocalMux I__6231 (
            .O(N__26286),
            .I(\ws2812.bit_counter_i_0 ));
    LocalMux I__6230 (
            .O(N__26283),
            .I(\ws2812.bit_counter_i_0 ));
    InMux I__6229 (
            .O(N__26278),
            .I(N__26275));
    LocalMux I__6228 (
            .O(N__26275),
            .I(\ws2812.un6_data_axb_1 ));
    InMux I__6227 (
            .O(N__26272),
            .I(\ws2812.un6_data_cry_0 ));
    InMux I__6226 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__6225 (
            .O(N__26266),
            .I(\ws2812.bit_counter_0_RNIQAT2Z0Z_0 ));
    InMux I__6224 (
            .O(N__26263),
            .I(\ws2812.un6_data_cry_1 ));
    InMux I__6223 (
            .O(N__26260),
            .I(N__26257));
    LocalMux I__6222 (
            .O(N__26257),
            .I(\ws2812.bit_counter_0_RNIRBT2Z0Z_1 ));
    InMux I__6221 (
            .O(N__26254),
            .I(\ws2812.un6_data_cry_2 ));
    InMux I__6220 (
            .O(N__26251),
            .I(N__26248));
    LocalMux I__6219 (
            .O(N__26248),
            .I(N__26245));
    Odrv4 I__6218 (
            .O(N__26245),
            .I(\ws2812.bit_counter_0_RNISCT2Z0Z_2 ));
    InMux I__6217 (
            .O(N__26242),
            .I(N__26236));
    InMux I__6216 (
            .O(N__26241),
            .I(N__26236));
    LocalMux I__6215 (
            .O(N__26236),
            .I(N__26233));
    Odrv4 I__6214 (
            .O(N__26233),
            .I(\ws2812.un6_data_cry_3_c_RNIKNFBZ0 ));
    InMux I__6213 (
            .O(N__26230),
            .I(\ws2812.un6_data_cry_3 ));
    InMux I__6212 (
            .O(N__26227),
            .I(N__26224));
    LocalMux I__6211 (
            .O(N__26224),
            .I(N__26221));
    Odrv4 I__6210 (
            .O(N__26221),
            .I(\ws2812.bit_counter_0_RNITDT2Z0Z_3 ));
    SRMux I__6209 (
            .O(N__26218),
            .I(N__26215));
    LocalMux I__6208 (
            .O(N__26215),
            .I(N__26204));
    SRMux I__6207 (
            .O(N__26214),
            .I(N__26201));
    SRMux I__6206 (
            .O(N__26213),
            .I(N__26198));
    SRMux I__6205 (
            .O(N__26212),
            .I(N__26192));
    CascadeMux I__6204 (
            .O(N__26211),
            .I(N__26188));
    CascadeMux I__6203 (
            .O(N__26210),
            .I(N__26185));
    CascadeMux I__6202 (
            .O(N__26209),
            .I(N__26182));
    CascadeMux I__6201 (
            .O(N__26208),
            .I(N__26179));
    SRMux I__6200 (
            .O(N__26207),
            .I(N__26174));
    Span4Mux_s2_v I__6199 (
            .O(N__26204),
            .I(N__26163));
    LocalMux I__6198 (
            .O(N__26201),
            .I(N__26163));
    LocalMux I__6197 (
            .O(N__26198),
            .I(N__26163));
    SRMux I__6196 (
            .O(N__26197),
            .I(N__26160));
    SRMux I__6195 (
            .O(N__26196),
            .I(N__26157));
    SRMux I__6194 (
            .O(N__26195),
            .I(N__26150));
    LocalMux I__6193 (
            .O(N__26192),
            .I(N__26145));
    SRMux I__6192 (
            .O(N__26191),
            .I(N__26142));
    InMux I__6191 (
            .O(N__26188),
            .I(N__26137));
    InMux I__6190 (
            .O(N__26185),
            .I(N__26137));
    InMux I__6189 (
            .O(N__26182),
            .I(N__26132));
    InMux I__6188 (
            .O(N__26179),
            .I(N__26132));
    SRMux I__6187 (
            .O(N__26178),
            .I(N__26129));
    SRMux I__6186 (
            .O(N__26177),
            .I(N__26126));
    LocalMux I__6185 (
            .O(N__26174),
            .I(N__26120));
    SRMux I__6184 (
            .O(N__26173),
            .I(N__26117));
    SRMux I__6183 (
            .O(N__26172),
            .I(N__26114));
    InMux I__6182 (
            .O(N__26171),
            .I(N__26111));
    SRMux I__6181 (
            .O(N__26170),
            .I(N__26108));
    Span4Mux_v I__6180 (
            .O(N__26163),
            .I(N__26101));
    LocalMux I__6179 (
            .O(N__26160),
            .I(N__26101));
    LocalMux I__6178 (
            .O(N__26157),
            .I(N__26101));
    SRMux I__6177 (
            .O(N__26156),
            .I(N__26098));
    SRMux I__6176 (
            .O(N__26155),
            .I(N__26094));
    SRMux I__6175 (
            .O(N__26154),
            .I(N__26091));
    SRMux I__6174 (
            .O(N__26153),
            .I(N__26088));
    LocalMux I__6173 (
            .O(N__26150),
            .I(N__26085));
    SRMux I__6172 (
            .O(N__26149),
            .I(N__26082));
    SRMux I__6171 (
            .O(N__26148),
            .I(N__26079));
    Span4Mux_v I__6170 (
            .O(N__26145),
            .I(N__26073));
    LocalMux I__6169 (
            .O(N__26142),
            .I(N__26073));
    LocalMux I__6168 (
            .O(N__26137),
            .I(N__26070));
    LocalMux I__6167 (
            .O(N__26132),
            .I(N__26067));
    LocalMux I__6166 (
            .O(N__26129),
            .I(N__26061));
    LocalMux I__6165 (
            .O(N__26126),
            .I(N__26061));
    SRMux I__6164 (
            .O(N__26125),
            .I(N__26058));
    DummyBuf I__6163 (
            .O(N__26124),
            .I(N__26055));
    DummyBuf I__6162 (
            .O(N__26123),
            .I(N__26052));
    Span4Mux_v I__6161 (
            .O(N__26120),
            .I(N__26045));
    LocalMux I__6160 (
            .O(N__26117),
            .I(N__26045));
    LocalMux I__6159 (
            .O(N__26114),
            .I(N__26045));
    LocalMux I__6158 (
            .O(N__26111),
            .I(N__26040));
    LocalMux I__6157 (
            .O(N__26108),
            .I(N__26040));
    Span4Mux_v I__6156 (
            .O(N__26101),
            .I(N__26035));
    LocalMux I__6155 (
            .O(N__26098),
            .I(N__26035));
    SRMux I__6154 (
            .O(N__26097),
            .I(N__26031));
    LocalMux I__6153 (
            .O(N__26094),
            .I(N__26028));
    LocalMux I__6152 (
            .O(N__26091),
            .I(N__26023));
    LocalMux I__6151 (
            .O(N__26088),
            .I(N__26023));
    Span4Mux_s1_v I__6150 (
            .O(N__26085),
            .I(N__26016));
    LocalMux I__6149 (
            .O(N__26082),
            .I(N__26016));
    LocalMux I__6148 (
            .O(N__26079),
            .I(N__26016));
    SRMux I__6147 (
            .O(N__26078),
            .I(N__26013));
    Span4Mux_v I__6146 (
            .O(N__26073),
            .I(N__26006));
    Span4Mux_s3_h I__6145 (
            .O(N__26070),
            .I(N__26006));
    Span4Mux_s3_h I__6144 (
            .O(N__26067),
            .I(N__26006));
    SRMux I__6143 (
            .O(N__26066),
            .I(N__26003));
    Span4Mux_v I__6142 (
            .O(N__26061),
            .I(N__25998));
    LocalMux I__6141 (
            .O(N__26058),
            .I(N__25998));
    InMux I__6140 (
            .O(N__26055),
            .I(N__25995));
    InMux I__6139 (
            .O(N__26052),
            .I(N__25992));
    Span4Mux_v I__6138 (
            .O(N__26045),
            .I(N__25985));
    Span4Mux_s3_h I__6137 (
            .O(N__26040),
            .I(N__25985));
    Span4Mux_s3_v I__6136 (
            .O(N__26035),
            .I(N__25985));
    SRMux I__6135 (
            .O(N__26034),
            .I(N__25982));
    LocalMux I__6134 (
            .O(N__26031),
            .I(N__25979));
    Span4Mux_h I__6133 (
            .O(N__26028),
            .I(N__25976));
    Span4Mux_v I__6132 (
            .O(N__26023),
            .I(N__25969));
    Span4Mux_v I__6131 (
            .O(N__26016),
            .I(N__25969));
    LocalMux I__6130 (
            .O(N__26013),
            .I(N__25969));
    Span4Mux_h I__6129 (
            .O(N__26006),
            .I(N__25964));
    LocalMux I__6128 (
            .O(N__26003),
            .I(N__25964));
    Span4Mux_h I__6127 (
            .O(N__25998),
            .I(N__25957));
    LocalMux I__6126 (
            .O(N__25995),
            .I(N__25957));
    LocalMux I__6125 (
            .O(N__25992),
            .I(N__25957));
    Span4Mux_h I__6124 (
            .O(N__25985),
            .I(N__25952));
    LocalMux I__6123 (
            .O(N__25982),
            .I(N__25952));
    Sp12to4 I__6122 (
            .O(N__25979),
            .I(N__25946));
    Span4Mux_h I__6121 (
            .O(N__25976),
            .I(N__25941));
    Span4Mux_v I__6120 (
            .O(N__25969),
            .I(N__25941));
    Span4Mux_h I__6119 (
            .O(N__25964),
            .I(N__25938));
    Span4Mux_v I__6118 (
            .O(N__25957),
            .I(N__25935));
    Span4Mux_h I__6117 (
            .O(N__25952),
            .I(N__25932));
    SRMux I__6116 (
            .O(N__25951),
            .I(N__25929));
    SRMux I__6115 (
            .O(N__25950),
            .I(N__25926));
    SRMux I__6114 (
            .O(N__25949),
            .I(N__25923));
    Odrv12 I__6113 (
            .O(N__25946),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6112 (
            .O(N__25941),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6111 (
            .O(N__25938),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6110 (
            .O(N__25935),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6109 (
            .O(N__25932),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6108 (
            .O(N__25929),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6107 (
            .O(N__25926),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6106 (
            .O(N__25923),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6105 (
            .O(N__25906),
            .I(N__25902));
    CascadeMux I__6104 (
            .O(N__25905),
            .I(N__25899));
    InMux I__6103 (
            .O(N__25902),
            .I(N__25894));
    InMux I__6102 (
            .O(N__25899),
            .I(N__25894));
    LocalMux I__6101 (
            .O(N__25894),
            .I(N__25891));
    Odrv4 I__6100 (
            .O(N__25891),
            .I(\ws2812.un6_data_cry_4_c_RNIMQGBZ0 ));
    InMux I__6099 (
            .O(N__25888),
            .I(\ws2812.un6_data_cry_4 ));
    InMux I__6098 (
            .O(N__25885),
            .I(N__25882));
    LocalMux I__6097 (
            .O(N__25882),
            .I(\ws2812.un6_data_axb_6 ));
    InMux I__6096 (
            .O(N__25879),
            .I(\ws2812.un6_data_cry_5 ));
    InMux I__6095 (
            .O(N__25876),
            .I(N__25873));
    LocalMux I__6094 (
            .O(N__25873),
            .I(\ws2812.un6_data_axb_7 ));
    InMux I__6093 (
            .O(N__25870),
            .I(\ws2812.un6_data_cry_6 ));
    CascadeMux I__6092 (
            .O(N__25867),
            .I(N__25863));
    InMux I__6091 (
            .O(N__25866),
            .I(N__25856));
    InMux I__6090 (
            .O(N__25863),
            .I(N__25845));
    InMux I__6089 (
            .O(N__25862),
            .I(N__25838));
    InMux I__6088 (
            .O(N__25861),
            .I(N__25838));
    InMux I__6087 (
            .O(N__25860),
            .I(N__25838));
    InMux I__6086 (
            .O(N__25859),
            .I(N__25833));
    LocalMux I__6085 (
            .O(N__25856),
            .I(N__25830));
    InMux I__6084 (
            .O(N__25855),
            .I(N__25821));
    InMux I__6083 (
            .O(N__25854),
            .I(N__25821));
    InMux I__6082 (
            .O(N__25853),
            .I(N__25821));
    InMux I__6081 (
            .O(N__25852),
            .I(N__25821));
    InMux I__6080 (
            .O(N__25851),
            .I(N__25816));
    InMux I__6079 (
            .O(N__25850),
            .I(N__25816));
    InMux I__6078 (
            .O(N__25849),
            .I(N__25811));
    InMux I__6077 (
            .O(N__25848),
            .I(N__25811));
    LocalMux I__6076 (
            .O(N__25845),
            .I(N__25808));
    LocalMux I__6075 (
            .O(N__25838),
            .I(N__25805));
    InMux I__6074 (
            .O(N__25837),
            .I(N__25802));
    InMux I__6073 (
            .O(N__25836),
            .I(N__25799));
    LocalMux I__6072 (
            .O(N__25833),
            .I(N__25792));
    Span4Mux_v I__6071 (
            .O(N__25830),
            .I(N__25792));
    LocalMux I__6070 (
            .O(N__25821),
            .I(N__25792));
    LocalMux I__6069 (
            .O(N__25816),
            .I(N__25789));
    LocalMux I__6068 (
            .O(N__25811),
            .I(N__25782));
    Span4Mux_v I__6067 (
            .O(N__25808),
            .I(N__25782));
    Span4Mux_v I__6066 (
            .O(N__25805),
            .I(N__25782));
    LocalMux I__6065 (
            .O(N__25802),
            .I(N__25777));
    LocalMux I__6064 (
            .O(N__25799),
            .I(N__25777));
    Span4Mux_h I__6063 (
            .O(N__25792),
            .I(N__25774));
    Odrv4 I__6062 (
            .O(N__25789),
            .I(\demux.N_424_i_0_o2Z0Z_0 ));
    Odrv4 I__6061 (
            .O(N__25782),
            .I(\demux.N_424_i_0_o2Z0Z_0 ));
    Odrv4 I__6060 (
            .O(N__25777),
            .I(\demux.N_424_i_0_o2Z0Z_0 ));
    Odrv4 I__6059 (
            .O(N__25774),
            .I(\demux.N_424_i_0_o2Z0Z_0 ));
    InMux I__6058 (
            .O(N__25765),
            .I(N__25761));
    InMux I__6057 (
            .O(N__25764),
            .I(N__25758));
    LocalMux I__6056 (
            .O(N__25761),
            .I(N__25754));
    LocalMux I__6055 (
            .O(N__25758),
            .I(N__25751));
    InMux I__6054 (
            .O(N__25757),
            .I(N__25748));
    Span4Mux_v I__6053 (
            .O(N__25754),
            .I(N__25744));
    Span4Mux_v I__6052 (
            .O(N__25751),
            .I(N__25739));
    LocalMux I__6051 (
            .O(N__25748),
            .I(N__25739));
    InMux I__6050 (
            .O(N__25747),
            .I(N__25736));
    Span4Mux_h I__6049 (
            .O(N__25744),
            .I(N__25733));
    Span4Mux_h I__6048 (
            .O(N__25739),
            .I(N__25728));
    LocalMux I__6047 (
            .O(N__25736),
            .I(N__25728));
    Odrv4 I__6046 (
            .O(N__25733),
            .I(\demux.N_419_i_0_o2Z0Z_9 ));
    Odrv4 I__6045 (
            .O(N__25728),
            .I(\demux.N_419_i_0_o2Z0Z_9 ));
    CascadeMux I__6044 (
            .O(N__25723),
            .I(N__25719));
    CascadeMux I__6043 (
            .O(N__25722),
            .I(N__25716));
    InMux I__6042 (
            .O(N__25719),
            .I(N__25712));
    InMux I__6041 (
            .O(N__25716),
            .I(N__25708));
    CascadeMux I__6040 (
            .O(N__25715),
            .I(N__25705));
    LocalMux I__6039 (
            .O(N__25712),
            .I(N__25702));
    CascadeMux I__6038 (
            .O(N__25711),
            .I(N__25699));
    LocalMux I__6037 (
            .O(N__25708),
            .I(N__25696));
    InMux I__6036 (
            .O(N__25705),
            .I(N__25693));
    Span4Mux_h I__6035 (
            .O(N__25702),
            .I(N__25690));
    InMux I__6034 (
            .O(N__25699),
            .I(N__25687));
    Span4Mux_s3_h I__6033 (
            .O(N__25696),
            .I(N__25682));
    LocalMux I__6032 (
            .O(N__25693),
            .I(N__25682));
    Sp12to4 I__6031 (
            .O(N__25690),
            .I(N__25677));
    LocalMux I__6030 (
            .O(N__25687),
            .I(N__25677));
    Span4Mux_v I__6029 (
            .O(N__25682),
            .I(N__25674));
    Span12Mux_v I__6028 (
            .O(N__25677),
            .I(N__25671));
    Sp12to4 I__6027 (
            .O(N__25674),
            .I(N__25668));
    Odrv12 I__6026 (
            .O(N__25671),
            .I(demux_data_in_5));
    Odrv12 I__6025 (
            .O(N__25668),
            .I(demux_data_in_5));
    InMux I__6024 (
            .O(N__25663),
            .I(N__25660));
    LocalMux I__6023 (
            .O(N__25660),
            .I(N__25657));
    Span4Mux_s2_h I__6022 (
            .O(N__25657),
            .I(N__25651));
    InMux I__6021 (
            .O(N__25656),
            .I(N__25648));
    InMux I__6020 (
            .O(N__25655),
            .I(N__25645));
    InMux I__6019 (
            .O(N__25654),
            .I(N__25642));
    Odrv4 I__6018 (
            .O(N__25651),
            .I(\demux.N_419_i_0_o2Z0Z_10 ));
    LocalMux I__6017 (
            .O(N__25648),
            .I(\demux.N_419_i_0_o2Z0Z_10 ));
    LocalMux I__6016 (
            .O(N__25645),
            .I(\demux.N_419_i_0_o2Z0Z_10 ));
    LocalMux I__6015 (
            .O(N__25642),
            .I(\demux.N_419_i_0_o2Z0Z_10 ));
    InMux I__6014 (
            .O(N__25633),
            .I(N__25630));
    LocalMux I__6013 (
            .O(N__25630),
            .I(N__25627));
    Odrv4 I__6012 (
            .O(N__25627),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_5 ));
    InMux I__6011 (
            .O(N__25624),
            .I(N__25619));
    InMux I__6010 (
            .O(N__25623),
            .I(N__25616));
    InMux I__6009 (
            .O(N__25622),
            .I(N__25613));
    LocalMux I__6008 (
            .O(N__25619),
            .I(N__25610));
    LocalMux I__6007 (
            .O(N__25616),
            .I(N__25607));
    LocalMux I__6006 (
            .O(N__25613),
            .I(N__25604));
    Span4Mux_s3_h I__6005 (
            .O(N__25610),
            .I(N__25600));
    Span4Mux_h I__6004 (
            .O(N__25607),
            .I(N__25597));
    Span4Mux_s3_h I__6003 (
            .O(N__25604),
            .I(N__25594));
    InMux I__6002 (
            .O(N__25603),
            .I(N__25591));
    Odrv4 I__6001 (
            .O(N__25600),
            .I(\demux.N_420_i_0_o2Z0Z_8 ));
    Odrv4 I__6000 (
            .O(N__25597),
            .I(\demux.N_420_i_0_o2Z0Z_8 ));
    Odrv4 I__5999 (
            .O(N__25594),
            .I(\demux.N_420_i_0_o2Z0Z_8 ));
    LocalMux I__5998 (
            .O(N__25591),
            .I(\demux.N_420_i_0_o2Z0Z_8 ));
    InMux I__5997 (
            .O(N__25582),
            .I(N__25578));
    InMux I__5996 (
            .O(N__25581),
            .I(N__25575));
    LocalMux I__5995 (
            .O(N__25578),
            .I(N__25571));
    LocalMux I__5994 (
            .O(N__25575),
            .I(N__25567));
    InMux I__5993 (
            .O(N__25574),
            .I(N__25564));
    Span4Mux_v I__5992 (
            .O(N__25571),
            .I(N__25561));
    InMux I__5991 (
            .O(N__25570),
            .I(N__25558));
    Span4Mux_v I__5990 (
            .O(N__25567),
            .I(N__25553));
    LocalMux I__5989 (
            .O(N__25564),
            .I(N__25553));
    Sp12to4 I__5988 (
            .O(N__25561),
            .I(N__25548));
    LocalMux I__5987 (
            .O(N__25558),
            .I(N__25548));
    Span4Mux_h I__5986 (
            .O(N__25553),
            .I(N__25545));
    Odrv12 I__5985 (
            .O(N__25548),
            .I(\demux.N_420_i_0_o2Z0Z_9 ));
    Odrv4 I__5984 (
            .O(N__25545),
            .I(\demux.N_420_i_0_o2Z0Z_9 ));
    CascadeMux I__5983 (
            .O(N__25540),
            .I(N__25535));
    CascadeMux I__5982 (
            .O(N__25539),
            .I(N__25531));
    CascadeMux I__5981 (
            .O(N__25538),
            .I(N__25528));
    InMux I__5980 (
            .O(N__25535),
            .I(N__25525));
    CascadeMux I__5979 (
            .O(N__25534),
            .I(N__25522));
    InMux I__5978 (
            .O(N__25531),
            .I(N__25519));
    InMux I__5977 (
            .O(N__25528),
            .I(N__25516));
    LocalMux I__5976 (
            .O(N__25525),
            .I(N__25513));
    InMux I__5975 (
            .O(N__25522),
            .I(N__25510));
    LocalMux I__5974 (
            .O(N__25519),
            .I(N__25507));
    LocalMux I__5973 (
            .O(N__25516),
            .I(N__25504));
    Span4Mux_v I__5972 (
            .O(N__25513),
            .I(N__25499));
    LocalMux I__5971 (
            .O(N__25510),
            .I(N__25499));
    Span4Mux_v I__5970 (
            .O(N__25507),
            .I(N__25494));
    Span4Mux_v I__5969 (
            .O(N__25504),
            .I(N__25494));
    Span4Mux_h I__5968 (
            .O(N__25499),
            .I(N__25491));
    Odrv4 I__5967 (
            .O(N__25494),
            .I(\demux.N_420_i_0_aZ0Z3 ));
    Odrv4 I__5966 (
            .O(N__25491),
            .I(\demux.N_420_i_0_aZ0Z3 ));
    InMux I__5965 (
            .O(N__25486),
            .I(N__25481));
    InMux I__5964 (
            .O(N__25485),
            .I(N__25478));
    InMux I__5963 (
            .O(N__25484),
            .I(N__25474));
    LocalMux I__5962 (
            .O(N__25481),
            .I(N__25471));
    LocalMux I__5961 (
            .O(N__25478),
            .I(N__25468));
    InMux I__5960 (
            .O(N__25477),
            .I(N__25465));
    LocalMux I__5959 (
            .O(N__25474),
            .I(N__25460));
    Span4Mux_s3_h I__5958 (
            .O(N__25471),
            .I(N__25460));
    Span4Mux_s3_h I__5957 (
            .O(N__25468),
            .I(N__25457));
    LocalMux I__5956 (
            .O(N__25465),
            .I(\demux.N_420_i_0_o2Z0Z_7 ));
    Odrv4 I__5955 (
            .O(N__25460),
            .I(\demux.N_420_i_0_o2Z0Z_7 ));
    Odrv4 I__5954 (
            .O(N__25457),
            .I(\demux.N_420_i_0_o2Z0Z_7 ));
    InMux I__5953 (
            .O(N__25450),
            .I(N__25447));
    LocalMux I__5952 (
            .O(N__25447),
            .I(N__25444));
    Odrv4 I__5951 (
            .O(N__25444),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_4 ));
    CEMux I__5950 (
            .O(N__25441),
            .I(N__25438));
    LocalMux I__5949 (
            .O(N__25438),
            .I(N__25434));
    CEMux I__5948 (
            .O(N__25437),
            .I(N__25431));
    Span4Mux_h I__5947 (
            .O(N__25434),
            .I(N__25425));
    LocalMux I__5946 (
            .O(N__25431),
            .I(N__25425));
    CEMux I__5945 (
            .O(N__25430),
            .I(N__25422));
    Span4Mux_v I__5944 (
            .O(N__25425),
            .I(N__25417));
    LocalMux I__5943 (
            .O(N__25422),
            .I(N__25417));
    Span4Mux_h I__5942 (
            .O(N__25417),
            .I(N__25414));
    Span4Mux_v I__5941 (
            .O(N__25414),
            .I(N__25411));
    Odrv4 I__5940 (
            .O(N__25411),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1 ));
    InMux I__5939 (
            .O(N__25408),
            .I(N__25404));
    InMux I__5938 (
            .O(N__25407),
            .I(N__25390));
    LocalMux I__5937 (
            .O(N__25404),
            .I(N__25387));
    InMux I__5936 (
            .O(N__25403),
            .I(N__25370));
    InMux I__5935 (
            .O(N__25402),
            .I(N__25370));
    InMux I__5934 (
            .O(N__25401),
            .I(N__25370));
    InMux I__5933 (
            .O(N__25400),
            .I(N__25370));
    InMux I__5932 (
            .O(N__25399),
            .I(N__25370));
    InMux I__5931 (
            .O(N__25398),
            .I(N__25370));
    InMux I__5930 (
            .O(N__25397),
            .I(N__25370));
    InMux I__5929 (
            .O(N__25396),
            .I(N__25370));
    CascadeMux I__5928 (
            .O(N__25395),
            .I(N__25366));
    CascadeMux I__5927 (
            .O(N__25394),
            .I(N__25362));
    CascadeMux I__5926 (
            .O(N__25393),
            .I(N__25357));
    LocalMux I__5925 (
            .O(N__25390),
            .I(N__25352));
    Span4Mux_v I__5924 (
            .O(N__25387),
            .I(N__25347));
    LocalMux I__5923 (
            .O(N__25370),
            .I(N__25347));
    InMux I__5922 (
            .O(N__25369),
            .I(N__25342));
    InMux I__5921 (
            .O(N__25366),
            .I(N__25342));
    InMux I__5920 (
            .O(N__25365),
            .I(N__25339));
    InMux I__5919 (
            .O(N__25362),
            .I(N__25326));
    InMux I__5918 (
            .O(N__25361),
            .I(N__25326));
    InMux I__5917 (
            .O(N__25360),
            .I(N__25326));
    InMux I__5916 (
            .O(N__25357),
            .I(N__25326));
    InMux I__5915 (
            .O(N__25356),
            .I(N__25326));
    InMux I__5914 (
            .O(N__25355),
            .I(N__25326));
    Span4Mux_v I__5913 (
            .O(N__25352),
            .I(N__25319));
    Span4Mux_h I__5912 (
            .O(N__25347),
            .I(N__25319));
    LocalMux I__5911 (
            .O(N__25342),
            .I(N__25319));
    LocalMux I__5910 (
            .O(N__25339),
            .I(\ws2812.stateZ0Z_1 ));
    LocalMux I__5909 (
            .O(N__25326),
            .I(\ws2812.stateZ0Z_1 ));
    Odrv4 I__5908 (
            .O(N__25319),
            .I(\ws2812.stateZ0Z_1 ));
    InMux I__5907 (
            .O(N__25312),
            .I(N__25306));
    InMux I__5906 (
            .O(N__25311),
            .I(N__25306));
    LocalMux I__5905 (
            .O(N__25306),
            .I(\ws2812.state_ns_0_i_o2_8_0 ));
    CascadeMux I__5904 (
            .O(N__25303),
            .I(N__25300));
    InMux I__5903 (
            .O(N__25300),
            .I(N__25297));
    LocalMux I__5902 (
            .O(N__25297),
            .I(N__25291));
    InMux I__5901 (
            .O(N__25296),
            .I(N__25288));
    InMux I__5900 (
            .O(N__25295),
            .I(N__25283));
    InMux I__5899 (
            .O(N__25294),
            .I(N__25283));
    Odrv12 I__5898 (
            .O(N__25291),
            .I(\ws2812.bit_counterZ0Z_1 ));
    LocalMux I__5897 (
            .O(N__25288),
            .I(\ws2812.bit_counterZ0Z_1 ));
    LocalMux I__5896 (
            .O(N__25283),
            .I(\ws2812.bit_counterZ0Z_1 ));
    InMux I__5895 (
            .O(N__25276),
            .I(N__25271));
    CascadeMux I__5894 (
            .O(N__25275),
            .I(N__25267));
    InMux I__5893 (
            .O(N__25274),
            .I(N__25264));
    LocalMux I__5892 (
            .O(N__25271),
            .I(N__25261));
    InMux I__5891 (
            .O(N__25270),
            .I(N__25258));
    InMux I__5890 (
            .O(N__25267),
            .I(N__25253));
    LocalMux I__5889 (
            .O(N__25264),
            .I(N__25248));
    Span4Mux_v I__5888 (
            .O(N__25261),
            .I(N__25248));
    LocalMux I__5887 (
            .O(N__25258),
            .I(N__25245));
    InMux I__5886 (
            .O(N__25257),
            .I(N__25240));
    InMux I__5885 (
            .O(N__25256),
            .I(N__25240));
    LocalMux I__5884 (
            .O(N__25253),
            .I(\ws2812.bit_counterZ0Z_0 ));
    Odrv4 I__5883 (
            .O(N__25248),
            .I(\ws2812.bit_counterZ0Z_0 ));
    Odrv4 I__5882 (
            .O(N__25245),
            .I(\ws2812.bit_counterZ0Z_0 ));
    LocalMux I__5881 (
            .O(N__25240),
            .I(\ws2812.bit_counterZ0Z_0 ));
    CascadeMux I__5880 (
            .O(N__25231),
            .I(N__25227));
    CascadeMux I__5879 (
            .O(N__25230),
            .I(N__25223));
    InMux I__5878 (
            .O(N__25227),
            .I(N__25220));
    InMux I__5877 (
            .O(N__25226),
            .I(N__25215));
    InMux I__5876 (
            .O(N__25223),
            .I(N__25215));
    LocalMux I__5875 (
            .O(N__25220),
            .I(N__25212));
    LocalMux I__5874 (
            .O(N__25215),
            .I(N__25209));
    Odrv4 I__5873 (
            .O(N__25212),
            .I(\ws2812.bit_counter_11 ));
    Odrv4 I__5872 (
            .O(N__25209),
            .I(\ws2812.bit_counter_11 ));
    InMux I__5871 (
            .O(N__25204),
            .I(N__25201));
    LocalMux I__5870 (
            .O(N__25201),
            .I(N__25198));
    Odrv4 I__5869 (
            .O(N__25198),
            .I(\ws2812.bit_counter_0_RNO_0Z0Z_4 ));
    InMux I__5868 (
            .O(N__25195),
            .I(N__25192));
    LocalMux I__5867 (
            .O(N__25192),
            .I(\ws2812.bit_counter_0_RNO_0Z0Z_0 ));
    CascadeMux I__5866 (
            .O(N__25189),
            .I(N__25186));
    InMux I__5865 (
            .O(N__25186),
            .I(N__25183));
    LocalMux I__5864 (
            .O(N__25183),
            .I(N__25177));
    InMux I__5863 (
            .O(N__25182),
            .I(N__25170));
    InMux I__5862 (
            .O(N__25181),
            .I(N__25170));
    InMux I__5861 (
            .O(N__25180),
            .I(N__25170));
    Odrv4 I__5860 (
            .O(N__25177),
            .I(\ws2812.bit_counterZ0Z_2 ));
    LocalMux I__5859 (
            .O(N__25170),
            .I(\ws2812.bit_counterZ0Z_2 ));
    InMux I__5858 (
            .O(N__25165),
            .I(N__25162));
    LocalMux I__5857 (
            .O(N__25162),
            .I(N__25159));
    Span4Mux_v I__5856 (
            .O(N__25159),
            .I(N__25156));
    Odrv4 I__5855 (
            .O(N__25156),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_13 ));
    InMux I__5854 (
            .O(N__25153),
            .I(N__25150));
    LocalMux I__5853 (
            .O(N__25150),
            .I(rgb_data_out_13));
    InMux I__5852 (
            .O(N__25147),
            .I(N__25144));
    LocalMux I__5851 (
            .O(N__25144),
            .I(N__25141));
    Span4Mux_h I__5850 (
            .O(N__25141),
            .I(N__25138));
    Odrv4 I__5849 (
            .O(N__25138),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_11 ));
    InMux I__5848 (
            .O(N__25135),
            .I(N__25132));
    LocalMux I__5847 (
            .O(N__25132),
            .I(N__25129));
    Odrv4 I__5846 (
            .O(N__25129),
            .I(rgb_data_out_11));
    InMux I__5845 (
            .O(N__25126),
            .I(N__25123));
    LocalMux I__5844 (
            .O(N__25123),
            .I(N__25120));
    Span4Mux_h I__5843 (
            .O(N__25120),
            .I(N__25117));
    Odrv4 I__5842 (
            .O(N__25117),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_9 ));
    InMux I__5841 (
            .O(N__25114),
            .I(N__25111));
    LocalMux I__5840 (
            .O(N__25111),
            .I(N__25108));
    Odrv4 I__5839 (
            .O(N__25108),
            .I(rgb_data_out_9));
    InMux I__5838 (
            .O(N__25105),
            .I(N__25102));
    LocalMux I__5837 (
            .O(N__25102),
            .I(N__25099));
    Odrv4 I__5836 (
            .O(N__25099),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_1 ));
    InMux I__5835 (
            .O(N__25096),
            .I(N__25093));
    LocalMux I__5834 (
            .O(N__25093),
            .I(N__25090));
    Span4Mux_s3_h I__5833 (
            .O(N__25090),
            .I(N__25087));
    Odrv4 I__5832 (
            .O(N__25087),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_21 ));
    InMux I__5831 (
            .O(N__25084),
            .I(N__25081));
    LocalMux I__5830 (
            .O(N__25081),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_20 ));
    CEMux I__5829 (
            .O(N__25078),
            .I(N__25074));
    CEMux I__5828 (
            .O(N__25077),
            .I(N__25071));
    LocalMux I__5827 (
            .O(N__25074),
            .I(N__25068));
    LocalMux I__5826 (
            .O(N__25071),
            .I(N__25065));
    Span4Mux_s3_h I__5825 (
            .O(N__25068),
            .I(N__25062));
    Span4Mux_v I__5824 (
            .O(N__25065),
            .I(N__25059));
    Span4Mux_v I__5823 (
            .O(N__25062),
            .I(N__25053));
    Span4Mux_s3_h I__5822 (
            .O(N__25059),
            .I(N__25053));
    CEMux I__5821 (
            .O(N__25058),
            .I(N__25050));
    Span4Mux_h I__5820 (
            .O(N__25053),
            .I(N__25047));
    LocalMux I__5819 (
            .O(N__25050),
            .I(N__25044));
    Odrv4 I__5818 (
            .O(N__25047),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1 ));
    Odrv12 I__5817 (
            .O(N__25044),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1 ));
    InMux I__5816 (
            .O(N__25039),
            .I(N__25036));
    LocalMux I__5815 (
            .O(N__25036),
            .I(N__25033));
    Span4Mux_s3_h I__5814 (
            .O(N__25033),
            .I(N__25030));
    Odrv4 I__5813 (
            .O(N__25030),
            .I(rgb_data_out_12));
    InMux I__5812 (
            .O(N__25027),
            .I(N__25024));
    LocalMux I__5811 (
            .O(N__25024),
            .I(N__25021));
    Span4Mux_s3_h I__5810 (
            .O(N__25021),
            .I(N__25018));
    Odrv4 I__5809 (
            .O(N__25018),
            .I(rgb_data_out_15));
    InMux I__5808 (
            .O(N__25015),
            .I(N__25012));
    LocalMux I__5807 (
            .O(N__25012),
            .I(N__25009));
    Span4Mux_s3_h I__5806 (
            .O(N__25009),
            .I(N__25006));
    Odrv4 I__5805 (
            .O(N__25006),
            .I(rgb_data_out_10));
    CascadeMux I__5804 (
            .O(N__25003),
            .I(\ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_ ));
    InMux I__5803 (
            .O(N__25000),
            .I(N__24997));
    LocalMux I__5802 (
            .O(N__24997),
            .I(\ws2812.rgb_counter_RNI2H7OZ0Z_2 ));
    InMux I__5801 (
            .O(N__24994),
            .I(N__24991));
    LocalMux I__5800 (
            .O(N__24991),
            .I(\ws2812.rgb_counter_RNIFI3MZ0Z_2 ));
    CascadeMux I__5799 (
            .O(N__24988),
            .I(\ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_ ));
    CascadeMux I__5798 (
            .O(N__24985),
            .I(\ws2812.N_108_cascade_ ));
    InMux I__5797 (
            .O(N__24982),
            .I(N__24976));
    InMux I__5796 (
            .O(N__24981),
            .I(N__24976));
    LocalMux I__5795 (
            .O(N__24976),
            .I(\ws2812.N_107 ));
    InMux I__5794 (
            .O(N__24973),
            .I(N__24970));
    LocalMux I__5793 (
            .O(N__24970),
            .I(\ws2812.rgb_counter_RNI4J7OZ0Z_2 ));
    InMux I__5792 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__5791 (
            .O(N__24964),
            .I(N__24961));
    Span4Mux_h I__5790 (
            .O(N__24961),
            .I(N__24958));
    Odrv4 I__5789 (
            .O(N__24958),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_8 ));
    InMux I__5788 (
            .O(N__24955),
            .I(N__24952));
    LocalMux I__5787 (
            .O(N__24952),
            .I(rgb_data_out_8));
    CascadeMux I__5786 (
            .O(N__24949),
            .I(N__24946));
    InMux I__5785 (
            .O(N__24946),
            .I(N__24943));
    LocalMux I__5784 (
            .O(N__24943),
            .I(N__24940));
    Odrv4 I__5783 (
            .O(N__24940),
            .I(\ws2812.bit_counter_RNI9RQB3Z0Z_5 ));
    InMux I__5782 (
            .O(N__24937),
            .I(\ws2812.un1_bit_counter_12_cry_8 ));
    CascadeMux I__5781 (
            .O(N__24934),
            .I(N__24931));
    InMux I__5780 (
            .O(N__24931),
            .I(N__24928));
    LocalMux I__5779 (
            .O(N__24928),
            .I(N__24925));
    Odrv12 I__5778 (
            .O(N__24925),
            .I(\ws2812.bit_counter_0_RNING643Z0Z_4 ));
    InMux I__5777 (
            .O(N__24922),
            .I(\ws2812.un1_bit_counter_12_cry_9 ));
    InMux I__5776 (
            .O(N__24919),
            .I(N__24916));
    LocalMux I__5775 (
            .O(N__24916),
            .I(N__24913));
    Odrv4 I__5774 (
            .O(N__24913),
            .I(\ws2812.un1_bit_counter_12_axb_11 ));
    InMux I__5773 (
            .O(N__24910),
            .I(\ws2812.un1_bit_counter_12_cry_10 ));
    InMux I__5772 (
            .O(N__24907),
            .I(N__24901));
    InMux I__5771 (
            .O(N__24906),
            .I(N__24901));
    LocalMux I__5770 (
            .O(N__24901),
            .I(N__24898));
    Odrv4 I__5769 (
            .O(N__24898),
            .I(\ws2812.state_ns_0_i_o2_7_0 ));
    InMux I__5768 (
            .O(N__24895),
            .I(N__24890));
    InMux I__5767 (
            .O(N__24894),
            .I(N__24884));
    InMux I__5766 (
            .O(N__24893),
            .I(N__24884));
    LocalMux I__5765 (
            .O(N__24890),
            .I(N__24881));
    InMux I__5764 (
            .O(N__24889),
            .I(N__24878));
    LocalMux I__5763 (
            .O(N__24884),
            .I(N__24875));
    Odrv12 I__5762 (
            .O(N__24881),
            .I(\ws2812.bit_counterZ0Z_4 ));
    LocalMux I__5761 (
            .O(N__24878),
            .I(\ws2812.bit_counterZ0Z_4 ));
    Odrv4 I__5760 (
            .O(N__24875),
            .I(\ws2812.bit_counterZ0Z_4 ));
    CascadeMux I__5759 (
            .O(N__24868),
            .I(N__24865));
    InMux I__5758 (
            .O(N__24865),
            .I(N__24860));
    InMux I__5757 (
            .O(N__24864),
            .I(N__24854));
    InMux I__5756 (
            .O(N__24863),
            .I(N__24854));
    LocalMux I__5755 (
            .O(N__24860),
            .I(N__24851));
    InMux I__5754 (
            .O(N__24859),
            .I(N__24848));
    LocalMux I__5753 (
            .O(N__24854),
            .I(N__24845));
    Odrv4 I__5752 (
            .O(N__24851),
            .I(\ws2812.bit_counterZ0Z_5 ));
    LocalMux I__5751 (
            .O(N__24848),
            .I(\ws2812.bit_counterZ0Z_5 ));
    Odrv4 I__5750 (
            .O(N__24845),
            .I(\ws2812.bit_counterZ0Z_5 ));
    InMux I__5749 (
            .O(N__24838),
            .I(N__24835));
    LocalMux I__5748 (
            .O(N__24835),
            .I(N__24829));
    InMux I__5747 (
            .O(N__24834),
            .I(N__24826));
    InMux I__5746 (
            .O(N__24833),
            .I(N__24821));
    InMux I__5745 (
            .O(N__24832),
            .I(N__24821));
    Odrv12 I__5744 (
            .O(N__24829),
            .I(\ws2812.bit_counter_8 ));
    LocalMux I__5743 (
            .O(N__24826),
            .I(\ws2812.bit_counter_8 ));
    LocalMux I__5742 (
            .O(N__24821),
            .I(\ws2812.bit_counter_8 ));
    CascadeMux I__5741 (
            .O(N__24814),
            .I(\ws2812.N_52_cascade_ ));
    IoInMux I__5740 (
            .O(N__24811),
            .I(N__24808));
    LocalMux I__5739 (
            .O(N__24808),
            .I(N__24805));
    Span4Mux_s3_v I__5738 (
            .O(N__24805),
            .I(N__24801));
    InMux I__5737 (
            .O(N__24804),
            .I(N__24798));
    Odrv4 I__5736 (
            .O(N__24801),
            .I(led));
    LocalMux I__5735 (
            .O(N__24798),
            .I(led));
    CascadeMux I__5734 (
            .O(N__24793),
            .I(N__24790));
    InMux I__5733 (
            .O(N__24790),
            .I(N__24787));
    LocalMux I__5732 (
            .O(N__24787),
            .I(N__24784));
    Odrv4 I__5731 (
            .O(N__24784),
            .I(\ws2812.bit_counter_RNI5NQB3Z0Z_1 ));
    InMux I__5730 (
            .O(N__24781),
            .I(\ws2812.un1_bit_counter_12_cry_0 ));
    InMux I__5729 (
            .O(N__24778),
            .I(N__24775));
    LocalMux I__5728 (
            .O(N__24775),
            .I(\ws2812.bit_counter_0_RNIJC643Z0Z_0 ));
    InMux I__5727 (
            .O(N__24772),
            .I(\ws2812.un1_bit_counter_12_cry_1 ));
    CascadeMux I__5726 (
            .O(N__24769),
            .I(N__24766));
    InMux I__5725 (
            .O(N__24766),
            .I(N__24761));
    InMux I__5724 (
            .O(N__24765),
            .I(N__24755));
    InMux I__5723 (
            .O(N__24764),
            .I(N__24755));
    LocalMux I__5722 (
            .O(N__24761),
            .I(N__24752));
    InMux I__5721 (
            .O(N__24760),
            .I(N__24749));
    LocalMux I__5720 (
            .O(N__24755),
            .I(N__24746));
    Span4Mux_v I__5719 (
            .O(N__24752),
            .I(N__24741));
    LocalMux I__5718 (
            .O(N__24749),
            .I(N__24741));
    Span4Mux_h I__5717 (
            .O(N__24746),
            .I(N__24738));
    Odrv4 I__5716 (
            .O(N__24741),
            .I(\ws2812.bit_counterZ0Z_3 ));
    Odrv4 I__5715 (
            .O(N__24738),
            .I(\ws2812.bit_counterZ0Z_3 ));
    CascadeMux I__5714 (
            .O(N__24733),
            .I(N__24730));
    InMux I__5713 (
            .O(N__24730),
            .I(N__24727));
    LocalMux I__5712 (
            .O(N__24727),
            .I(N__24724));
    Odrv4 I__5711 (
            .O(N__24724),
            .I(\ws2812.bit_counter_0_RNIKD643Z0Z_1 ));
    InMux I__5710 (
            .O(N__24721),
            .I(N__24718));
    LocalMux I__5709 (
            .O(N__24718),
            .I(N__24715));
    Odrv4 I__5708 (
            .O(N__24715),
            .I(\ws2812.bit_counter_0_RNO_0Z0Z_1 ));
    InMux I__5707 (
            .O(N__24712),
            .I(\ws2812.un1_bit_counter_12_cry_2 ));
    CascadeMux I__5706 (
            .O(N__24709),
            .I(N__24706));
    InMux I__5705 (
            .O(N__24706),
            .I(N__24703));
    LocalMux I__5704 (
            .O(N__24703),
            .I(N__24700));
    Odrv4 I__5703 (
            .O(N__24700),
            .I(\ws2812.bit_counter_0_RNILE643Z0Z_2 ));
    InMux I__5702 (
            .O(N__24697),
            .I(\ws2812.un1_bit_counter_12_cry_3 ));
    CascadeMux I__5701 (
            .O(N__24694),
            .I(N__24691));
    InMux I__5700 (
            .O(N__24691),
            .I(N__24688));
    LocalMux I__5699 (
            .O(N__24688),
            .I(N__24685));
    Odrv4 I__5698 (
            .O(N__24685),
            .I(\ws2812.bit_counter_0_RNIMF643Z0Z_3 ));
    InMux I__5697 (
            .O(N__24682),
            .I(\ws2812.un1_bit_counter_12_cry_4 ));
    CascadeMux I__5696 (
            .O(N__24679),
            .I(N__24676));
    InMux I__5695 (
            .O(N__24676),
            .I(N__24673));
    LocalMux I__5694 (
            .O(N__24673),
            .I(N__24670));
    Span4Mux_h I__5693 (
            .O(N__24670),
            .I(N__24667));
    Odrv4 I__5692 (
            .O(N__24667),
            .I(\ws2812.bit_counter_RNI6OQB3Z0Z_2 ));
    InMux I__5691 (
            .O(N__24664),
            .I(N__24661));
    LocalMux I__5690 (
            .O(N__24661),
            .I(N__24658));
    Span12Mux_s9_v I__5689 (
            .O(N__24658),
            .I(N__24652));
    InMux I__5688 (
            .O(N__24657),
            .I(N__24649));
    InMux I__5687 (
            .O(N__24656),
            .I(N__24644));
    InMux I__5686 (
            .O(N__24655),
            .I(N__24644));
    Odrv12 I__5685 (
            .O(N__24652),
            .I(\ws2812.bit_counter_6 ));
    LocalMux I__5684 (
            .O(N__24649),
            .I(\ws2812.bit_counter_6 ));
    LocalMux I__5683 (
            .O(N__24644),
            .I(\ws2812.bit_counter_6 ));
    InMux I__5682 (
            .O(N__24637),
            .I(\ws2812.un1_bit_counter_12_cry_5 ));
    CascadeMux I__5681 (
            .O(N__24634),
            .I(N__24631));
    InMux I__5680 (
            .O(N__24631),
            .I(N__24628));
    LocalMux I__5679 (
            .O(N__24628),
            .I(N__24625));
    Span4Mux_s3_h I__5678 (
            .O(N__24625),
            .I(N__24622));
    Odrv4 I__5677 (
            .O(N__24622),
            .I(\ws2812.bit_counter_RNI7PQB3Z0Z_3 ));
    CascadeMux I__5676 (
            .O(N__24619),
            .I(N__24616));
    InMux I__5675 (
            .O(N__24616),
            .I(N__24613));
    LocalMux I__5674 (
            .O(N__24613),
            .I(N__24609));
    CascadeMux I__5673 (
            .O(N__24612),
            .I(N__24604));
    Span4Mux_v I__5672 (
            .O(N__24609),
            .I(N__24601));
    InMux I__5671 (
            .O(N__24608),
            .I(N__24598));
    InMux I__5670 (
            .O(N__24607),
            .I(N__24593));
    InMux I__5669 (
            .O(N__24604),
            .I(N__24593));
    Odrv4 I__5668 (
            .O(N__24601),
            .I(\ws2812.bit_counter_7 ));
    LocalMux I__5667 (
            .O(N__24598),
            .I(\ws2812.bit_counter_7 ));
    LocalMux I__5666 (
            .O(N__24593),
            .I(\ws2812.bit_counter_7 ));
    InMux I__5665 (
            .O(N__24586),
            .I(\ws2812.un1_bit_counter_12_cry_6 ));
    CascadeMux I__5664 (
            .O(N__24583),
            .I(N__24580));
    InMux I__5663 (
            .O(N__24580),
            .I(N__24577));
    LocalMux I__5662 (
            .O(N__24577),
            .I(N__24574));
    Odrv4 I__5661 (
            .O(N__24574),
            .I(\ws2812.bit_counter_RNI8QQB3Z0Z_4 ));
    InMux I__5660 (
            .O(N__24571),
            .I(bfn_11_6_0_));
    CascadeMux I__5659 (
            .O(N__24568),
            .I(\ws2812.state_ns_0_i_o2_6_0_cascade_ ));
    CascadeMux I__5658 (
            .O(N__24565),
            .I(\ws2812.N_105_cascade_ ));
    InMux I__5657 (
            .O(N__24562),
            .I(N__24559));
    LocalMux I__5656 (
            .O(N__24559),
            .I(\ws2812.state_ns_0_i_o2_6_0 ));
    CascadeMux I__5655 (
            .O(N__24556),
            .I(N__24553));
    InMux I__5654 (
            .O(N__24553),
            .I(N__24550));
    LocalMux I__5653 (
            .O(N__24550),
            .I(N__24547));
    Odrv4 I__5652 (
            .O(N__24547),
            .I(\ws2812.un1_bit_counter_12_cry_0_c_RNOZ0 ));
    InMux I__5651 (
            .O(N__24544),
            .I(N__24541));
    LocalMux I__5650 (
            .O(N__24541),
            .I(N__24538));
    Span4Mux_v I__5649 (
            .O(N__24538),
            .I(N__24535));
    Odrv4 I__5648 (
            .O(N__24535),
            .I(demux_data_in_101));
    InMux I__5647 (
            .O(N__24532),
            .I(N__24529));
    LocalMux I__5646 (
            .O(N__24529),
            .I(demux_data_in_21));
    InMux I__5645 (
            .O(N__24526),
            .I(N__24523));
    LocalMux I__5644 (
            .O(N__24523),
            .I(\demux.N_419_i_0_o2Z0Z_4 ));
    InMux I__5643 (
            .O(N__24520),
            .I(N__24517));
    LocalMux I__5642 (
            .O(N__24517),
            .I(N__24514));
    Span4Mux_v I__5641 (
            .O(N__24514),
            .I(N__24511));
    Odrv4 I__5640 (
            .O(N__24511),
            .I(demux_data_in_100));
    CascadeMux I__5639 (
            .O(N__24508),
            .I(N__24499));
    CascadeMux I__5638 (
            .O(N__24507),
            .I(N__24496));
    InMux I__5637 (
            .O(N__24506),
            .I(N__24493));
    InMux I__5636 (
            .O(N__24505),
            .I(N__24488));
    InMux I__5635 (
            .O(N__24504),
            .I(N__24488));
    InMux I__5634 (
            .O(N__24503),
            .I(N__24479));
    InMux I__5633 (
            .O(N__24502),
            .I(N__24479));
    InMux I__5632 (
            .O(N__24499),
            .I(N__24479));
    InMux I__5631 (
            .O(N__24496),
            .I(N__24479));
    LocalMux I__5630 (
            .O(N__24493),
            .I(N__24475));
    LocalMux I__5629 (
            .O(N__24488),
            .I(N__24472));
    LocalMux I__5628 (
            .O(N__24479),
            .I(N__24469));
    InMux I__5627 (
            .O(N__24478),
            .I(N__24466));
    Span4Mux_h I__5626 (
            .O(N__24475),
            .I(N__24463));
    Span4Mux_h I__5625 (
            .O(N__24472),
            .I(N__24458));
    Span4Mux_h I__5624 (
            .O(N__24469),
            .I(N__24458));
    LocalMux I__5623 (
            .O(N__24466),
            .I(\demux.N_424_i_0_a2Z0Z_3 ));
    Odrv4 I__5622 (
            .O(N__24463),
            .I(\demux.N_424_i_0_a2Z0Z_3 ));
    Odrv4 I__5621 (
            .O(N__24458),
            .I(\demux.N_424_i_0_a2Z0Z_3 ));
    CascadeMux I__5620 (
            .O(N__24451),
            .I(N__24448));
    InMux I__5619 (
            .O(N__24448),
            .I(N__24445));
    LocalMux I__5618 (
            .O(N__24445),
            .I(N__24442));
    Span4Mux_h I__5617 (
            .O(N__24442),
            .I(N__24439));
    Odrv4 I__5616 (
            .O(N__24439),
            .I(demux_data_in_20));
    InMux I__5615 (
            .O(N__24436),
            .I(N__24427));
    InMux I__5614 (
            .O(N__24435),
            .I(N__24424));
    InMux I__5613 (
            .O(N__24434),
            .I(N__24421));
    InMux I__5612 (
            .O(N__24433),
            .I(N__24412));
    InMux I__5611 (
            .O(N__24432),
            .I(N__24412));
    InMux I__5610 (
            .O(N__24431),
            .I(N__24412));
    InMux I__5609 (
            .O(N__24430),
            .I(N__24412));
    LocalMux I__5608 (
            .O(N__24427),
            .I(N__24408));
    LocalMux I__5607 (
            .O(N__24424),
            .I(N__24405));
    LocalMux I__5606 (
            .O(N__24421),
            .I(N__24402));
    LocalMux I__5605 (
            .O(N__24412),
            .I(N__24399));
    InMux I__5604 (
            .O(N__24411),
            .I(N__24396));
    Span4Mux_h I__5603 (
            .O(N__24408),
            .I(N__24393));
    Span4Mux_h I__5602 (
            .O(N__24405),
            .I(N__24390));
    Span4Mux_h I__5601 (
            .O(N__24402),
            .I(N__24385));
    Span4Mux_h I__5600 (
            .O(N__24399),
            .I(N__24385));
    LocalMux I__5599 (
            .O(N__24396),
            .I(\demux.N_424_i_0_a2Z0Z_10 ));
    Odrv4 I__5598 (
            .O(N__24393),
            .I(\demux.N_424_i_0_a2Z0Z_10 ));
    Odrv4 I__5597 (
            .O(N__24390),
            .I(\demux.N_424_i_0_a2Z0Z_10 ));
    Odrv4 I__5596 (
            .O(N__24385),
            .I(\demux.N_424_i_0_a2Z0Z_10 ));
    InMux I__5595 (
            .O(N__24376),
            .I(N__24373));
    LocalMux I__5594 (
            .O(N__24373),
            .I(N__24370));
    Span4Mux_h I__5593 (
            .O(N__24370),
            .I(N__24367));
    Span4Mux_h I__5592 (
            .O(N__24367),
            .I(N__24364));
    Odrv4 I__5591 (
            .O(N__24364),
            .I(demux_data_in_68));
    InMux I__5590 (
            .O(N__24361),
            .I(N__24355));
    CascadeMux I__5589 (
            .O(N__24360),
            .I(N__24350));
    InMux I__5588 (
            .O(N__24359),
            .I(N__24344));
    InMux I__5587 (
            .O(N__24358),
            .I(N__24344));
    LocalMux I__5586 (
            .O(N__24355),
            .I(N__24341));
    InMux I__5585 (
            .O(N__24354),
            .I(N__24338));
    InMux I__5584 (
            .O(N__24353),
            .I(N__24335));
    InMux I__5583 (
            .O(N__24350),
            .I(N__24330));
    InMux I__5582 (
            .O(N__24349),
            .I(N__24330));
    LocalMux I__5581 (
            .O(N__24344),
            .I(N__24327));
    Span4Mux_h I__5580 (
            .O(N__24341),
            .I(N__24321));
    LocalMux I__5579 (
            .O(N__24338),
            .I(N__24321));
    LocalMux I__5578 (
            .O(N__24335),
            .I(N__24318));
    LocalMux I__5577 (
            .O(N__24330),
            .I(N__24315));
    Span4Mux_s3_v I__5576 (
            .O(N__24327),
            .I(N__24312));
    InMux I__5575 (
            .O(N__24326),
            .I(N__24309));
    Span4Mux_v I__5574 (
            .O(N__24321),
            .I(N__24304));
    Span4Mux_s3_v I__5573 (
            .O(N__24318),
            .I(N__24304));
    Span4Mux_h I__5572 (
            .O(N__24315),
            .I(N__24301));
    Odrv4 I__5571 (
            .O(N__24312),
            .I(\demux.N_424_i_0_a2Z0Z_9 ));
    LocalMux I__5570 (
            .O(N__24309),
            .I(\demux.N_424_i_0_a2Z0Z_9 ));
    Odrv4 I__5569 (
            .O(N__24304),
            .I(\demux.N_424_i_0_a2Z0Z_9 ));
    Odrv4 I__5568 (
            .O(N__24301),
            .I(\demux.N_424_i_0_a2Z0Z_9 ));
    CascadeMux I__5567 (
            .O(N__24292),
            .I(\demux.N_420_i_0_o2Z0Z_4_cascade_ ));
    InMux I__5566 (
            .O(N__24289),
            .I(N__24286));
    LocalMux I__5565 (
            .O(N__24286),
            .I(N__24283));
    Span4Mux_h I__5564 (
            .O(N__24283),
            .I(N__24280));
    Odrv4 I__5563 (
            .O(N__24280),
            .I(\demux.N_420_i_0_a3Z0Z_7 ));
    InMux I__5562 (
            .O(N__24277),
            .I(N__24274));
    LocalMux I__5561 (
            .O(N__24274),
            .I(N__24271));
    Span12Mux_s9_h I__5560 (
            .O(N__24271),
            .I(N__24268));
    Odrv12 I__5559 (
            .O(N__24268),
            .I(miso_data_in_5));
    InMux I__5558 (
            .O(N__24265),
            .I(N__24260));
    InMux I__5557 (
            .O(N__24264),
            .I(N__24257));
    CascadeMux I__5556 (
            .O(N__24263),
            .I(N__24253));
    LocalMux I__5555 (
            .O(N__24260),
            .I(N__24248));
    LocalMux I__5554 (
            .O(N__24257),
            .I(N__24248));
    InMux I__5553 (
            .O(N__24256),
            .I(N__24245));
    InMux I__5552 (
            .O(N__24253),
            .I(N__24242));
    Span4Mux_v I__5551 (
            .O(N__24248),
            .I(N__24239));
    LocalMux I__5550 (
            .O(N__24245),
            .I(N__24236));
    LocalMux I__5549 (
            .O(N__24242),
            .I(N__24233));
    Span4Mux_h I__5548 (
            .O(N__24239),
            .I(N__24230));
    Span4Mux_h I__5547 (
            .O(N__24236),
            .I(N__24225));
    Span4Mux_v I__5546 (
            .O(N__24233),
            .I(N__24225));
    Odrv4 I__5545 (
            .O(N__24230),
            .I(\demux.N_421_i_0_o2Z0Z_9 ));
    Odrv4 I__5544 (
            .O(N__24225),
            .I(\demux.N_421_i_0_o2Z0Z_9 ));
    InMux I__5543 (
            .O(N__24220),
            .I(N__24215));
    InMux I__5542 (
            .O(N__24219),
            .I(N__24212));
    CascadeMux I__5541 (
            .O(N__24218),
            .I(N__24208));
    LocalMux I__5540 (
            .O(N__24215),
            .I(N__24205));
    LocalMux I__5539 (
            .O(N__24212),
            .I(N__24202));
    InMux I__5538 (
            .O(N__24211),
            .I(N__24199));
    InMux I__5537 (
            .O(N__24208),
            .I(N__24196));
    Span4Mux_h I__5536 (
            .O(N__24205),
            .I(N__24187));
    Span4Mux_v I__5535 (
            .O(N__24202),
            .I(N__24187));
    LocalMux I__5534 (
            .O(N__24199),
            .I(N__24187));
    LocalMux I__5533 (
            .O(N__24196),
            .I(N__24187));
    Span4Mux_v I__5532 (
            .O(N__24187),
            .I(N__24184));
    Span4Mux_v I__5531 (
            .O(N__24184),
            .I(N__24181));
    Odrv4 I__5530 (
            .O(N__24181),
            .I(demux_data_in_3));
    CascadeMux I__5529 (
            .O(N__24178),
            .I(N__24173));
    InMux I__5528 (
            .O(N__24177),
            .I(N__24169));
    InMux I__5527 (
            .O(N__24176),
            .I(N__24166));
    InMux I__5526 (
            .O(N__24173),
            .I(N__24163));
    InMux I__5525 (
            .O(N__24172),
            .I(N__24160));
    LocalMux I__5524 (
            .O(N__24169),
            .I(N__24157));
    LocalMux I__5523 (
            .O(N__24166),
            .I(N__24152));
    LocalMux I__5522 (
            .O(N__24163),
            .I(N__24152));
    LocalMux I__5521 (
            .O(N__24160),
            .I(\demux.N_421_i_0_o2Z0Z_10 ));
    Odrv4 I__5520 (
            .O(N__24157),
            .I(\demux.N_421_i_0_o2Z0Z_10 ));
    Odrv4 I__5519 (
            .O(N__24152),
            .I(\demux.N_421_i_0_o2Z0Z_10 ));
    InMux I__5518 (
            .O(N__24145),
            .I(N__24142));
    LocalMux I__5517 (
            .O(N__24142),
            .I(N__24139));
    Odrv12 I__5516 (
            .O(N__24139),
            .I(miso_data_in_3));
    CascadeMux I__5515 (
            .O(N__24136),
            .I(N__24132));
    InMux I__5514 (
            .O(N__24135),
            .I(N__24128));
    InMux I__5513 (
            .O(N__24132),
            .I(N__24125));
    InMux I__5512 (
            .O(N__24131),
            .I(N__24122));
    LocalMux I__5511 (
            .O(N__24128),
            .I(N__24118));
    LocalMux I__5510 (
            .O(N__24125),
            .I(N__24113));
    LocalMux I__5509 (
            .O(N__24122),
            .I(N__24113));
    InMux I__5508 (
            .O(N__24121),
            .I(N__24110));
    Span4Mux_v I__5507 (
            .O(N__24118),
            .I(N__24103));
    Span4Mux_v I__5506 (
            .O(N__24113),
            .I(N__24103));
    LocalMux I__5505 (
            .O(N__24110),
            .I(N__24103));
    Span4Mux_h I__5504 (
            .O(N__24103),
            .I(N__24100));
    Odrv4 I__5503 (
            .O(N__24100),
            .I(\demux.N_423_i_0_o2Z0Z_9 ));
    CascadeMux I__5502 (
            .O(N__24097),
            .I(N__24094));
    InMux I__5501 (
            .O(N__24094),
            .I(N__24089));
    InMux I__5500 (
            .O(N__24093),
            .I(N__24086));
    InMux I__5499 (
            .O(N__24092),
            .I(N__24082));
    LocalMux I__5498 (
            .O(N__24089),
            .I(N__24077));
    LocalMux I__5497 (
            .O(N__24086),
            .I(N__24077));
    CascadeMux I__5496 (
            .O(N__24085),
            .I(N__24074));
    LocalMux I__5495 (
            .O(N__24082),
            .I(N__24071));
    Span4Mux_v I__5494 (
            .O(N__24077),
            .I(N__24068));
    InMux I__5493 (
            .O(N__24074),
            .I(N__24065));
    Span4Mux_v I__5492 (
            .O(N__24071),
            .I(N__24062));
    Span4Mux_h I__5491 (
            .O(N__24068),
            .I(N__24057));
    LocalMux I__5490 (
            .O(N__24065),
            .I(N__24057));
    Span4Mux_v I__5489 (
            .O(N__24062),
            .I(N__24054));
    Span4Mux_v I__5488 (
            .O(N__24057),
            .I(N__24051));
    Odrv4 I__5487 (
            .O(N__24054),
            .I(demux_data_in_1));
    Odrv4 I__5486 (
            .O(N__24051),
            .I(demux_data_in_1));
    InMux I__5485 (
            .O(N__24046),
            .I(N__24040));
    InMux I__5484 (
            .O(N__24045),
            .I(N__24037));
    InMux I__5483 (
            .O(N__24044),
            .I(N__24034));
    InMux I__5482 (
            .O(N__24043),
            .I(N__24031));
    LocalMux I__5481 (
            .O(N__24040),
            .I(\demux.N_423_i_0_o2Z0Z_10 ));
    LocalMux I__5480 (
            .O(N__24037),
            .I(\demux.N_423_i_0_o2Z0Z_10 ));
    LocalMux I__5479 (
            .O(N__24034),
            .I(\demux.N_423_i_0_o2Z0Z_10 ));
    LocalMux I__5478 (
            .O(N__24031),
            .I(\demux.N_423_i_0_o2Z0Z_10 ));
    InMux I__5477 (
            .O(N__24022),
            .I(N__24019));
    LocalMux I__5476 (
            .O(N__24019),
            .I(N__24016));
    Odrv12 I__5475 (
            .O(N__24016),
            .I(miso_data_in_1));
    InMux I__5474 (
            .O(N__24013),
            .I(N__24010));
    LocalMux I__5473 (
            .O(N__24010),
            .I(N__24007));
    Span4Mux_h I__5472 (
            .O(N__24007),
            .I(N__24004));
    Span4Mux_h I__5471 (
            .O(N__24004),
            .I(N__24001));
    Odrv4 I__5470 (
            .O(N__24001),
            .I(miso_data_in_4));
    InMux I__5469 (
            .O(N__23998),
            .I(N__23995));
    LocalMux I__5468 (
            .O(N__23995),
            .I(N__23988));
    CEMux I__5467 (
            .O(N__23994),
            .I(N__23977));
    CEMux I__5466 (
            .O(N__23993),
            .I(N__23977));
    CEMux I__5465 (
            .O(N__23992),
            .I(N__23977));
    CEMux I__5464 (
            .O(N__23991),
            .I(N__23977));
    Glb2LocalMux I__5463 (
            .O(N__23988),
            .I(N__23977));
    GlobalMux I__5462 (
            .O(N__23977),
            .I(N__23974));
    gio2CtrlBuf I__5461 (
            .O(N__23974),
            .I(\sb_translator_1.state_g_1 ));
    InMux I__5460 (
            .O(N__23971),
            .I(N__23968));
    LocalMux I__5459 (
            .O(N__23968),
            .I(N__23965));
    Sp12to4 I__5458 (
            .O(N__23965),
            .I(N__23962));
    Span12Mux_v I__5457 (
            .O(N__23962),
            .I(N__23959));
    Odrv12 I__5456 (
            .O(N__23959),
            .I(demux_data_in_31));
    InMux I__5455 (
            .O(N__23956),
            .I(N__23952));
    InMux I__5454 (
            .O(N__23955),
            .I(N__23946));
    LocalMux I__5453 (
            .O(N__23952),
            .I(N__23943));
    InMux I__5452 (
            .O(N__23951),
            .I(N__23940));
    InMux I__5451 (
            .O(N__23950),
            .I(N__23935));
    InMux I__5450 (
            .O(N__23949),
            .I(N__23935));
    LocalMux I__5449 (
            .O(N__23946),
            .I(N__23932));
    Span4Mux_h I__5448 (
            .O(N__23943),
            .I(N__23923));
    LocalMux I__5447 (
            .O(N__23940),
            .I(N__23923));
    LocalMux I__5446 (
            .O(N__23935),
            .I(N__23923));
    Span4Mux_h I__5445 (
            .O(N__23932),
            .I(N__23919));
    InMux I__5444 (
            .O(N__23931),
            .I(N__23914));
    InMux I__5443 (
            .O(N__23930),
            .I(N__23914));
    Span4Mux_v I__5442 (
            .O(N__23923),
            .I(N__23911));
    InMux I__5441 (
            .O(N__23922),
            .I(N__23908));
    Odrv4 I__5440 (
            .O(N__23919),
            .I(\demux.N_424_i_0_a2Z0Z_1 ));
    LocalMux I__5439 (
            .O(N__23914),
            .I(\demux.N_424_i_0_a2Z0Z_1 ));
    Odrv4 I__5438 (
            .O(N__23911),
            .I(\demux.N_424_i_0_a2Z0Z_1 ));
    LocalMux I__5437 (
            .O(N__23908),
            .I(\demux.N_424_i_0_a2Z0Z_1 ));
    InMux I__5436 (
            .O(N__23899),
            .I(N__23896));
    LocalMux I__5435 (
            .O(N__23896),
            .I(N__23893));
    Span12Mux_s10_h I__5434 (
            .O(N__23893),
            .I(N__23890));
    Odrv12 I__5433 (
            .O(N__23890),
            .I(demux_data_in_71));
    CascadeMux I__5432 (
            .O(N__23887),
            .I(\demux.N_417_i_0_a3Z0Z_7_cascade_ ));
    InMux I__5431 (
            .O(N__23884),
            .I(N__23878));
    InMux I__5430 (
            .O(N__23883),
            .I(N__23875));
    InMux I__5429 (
            .O(N__23882),
            .I(N__23872));
    InMux I__5428 (
            .O(N__23881),
            .I(N__23869));
    LocalMux I__5427 (
            .O(N__23878),
            .I(N__23860));
    LocalMux I__5426 (
            .O(N__23875),
            .I(N__23860));
    LocalMux I__5425 (
            .O(N__23872),
            .I(N__23860));
    LocalMux I__5424 (
            .O(N__23869),
            .I(N__23860));
    Odrv4 I__5423 (
            .O(N__23860),
            .I(\demux.N_417_i_0_o2Z0Z_8 ));
    InMux I__5422 (
            .O(N__23857),
            .I(N__23854));
    LocalMux I__5421 (
            .O(N__23854),
            .I(N__23851));
    Span4Mux_v I__5420 (
            .O(N__23851),
            .I(N__23848));
    Odrv4 I__5419 (
            .O(N__23848),
            .I(demux_data_in_103));
    InMux I__5418 (
            .O(N__23845),
            .I(N__23842));
    LocalMux I__5417 (
            .O(N__23842),
            .I(demux_data_in_23));
    InMux I__5416 (
            .O(N__23839),
            .I(N__23836));
    LocalMux I__5415 (
            .O(N__23836),
            .I(\demux.N_417_i_0_o2Z0Z_4 ));
    InMux I__5414 (
            .O(N__23833),
            .I(N__23830));
    LocalMux I__5413 (
            .O(N__23830),
            .I(N__23827));
    Odrv4 I__5412 (
            .O(N__23827),
            .I(demux_data_in_18));
    CascadeMux I__5411 (
            .O(N__23824),
            .I(N__23821));
    InMux I__5410 (
            .O(N__23821),
            .I(N__23818));
    LocalMux I__5409 (
            .O(N__23818),
            .I(N__23815));
    Sp12to4 I__5408 (
            .O(N__23815),
            .I(N__23812));
    Odrv12 I__5407 (
            .O(N__23812),
            .I(demux_data_in_98));
    InMux I__5406 (
            .O(N__23809),
            .I(N__23806));
    LocalMux I__5405 (
            .O(N__23806),
            .I(N__23803));
    Span4Mux_v I__5404 (
            .O(N__23803),
            .I(N__23800));
    Odrv4 I__5403 (
            .O(N__23800),
            .I(\demux.N_422_i_0_o2Z0Z_4 ));
    CascadeMux I__5402 (
            .O(N__23797),
            .I(\demux.N_874_cascade_ ));
    InMux I__5401 (
            .O(N__23794),
            .I(N__23791));
    LocalMux I__5400 (
            .O(N__23791),
            .I(N__23788));
    Span4Mux_v I__5399 (
            .O(N__23788),
            .I(N__23785));
    Span4Mux_v I__5398 (
            .O(N__23785),
            .I(N__23782));
    Odrv4 I__5397 (
            .O(N__23782),
            .I(demux_data_in_4));
    InMux I__5396 (
            .O(N__23779),
            .I(N__23775));
    InMux I__5395 (
            .O(N__23778),
            .I(N__23772));
    LocalMux I__5394 (
            .O(N__23775),
            .I(N__23767));
    LocalMux I__5393 (
            .O(N__23772),
            .I(N__23764));
    InMux I__5392 (
            .O(N__23771),
            .I(N__23761));
    InMux I__5391 (
            .O(N__23770),
            .I(N__23758));
    Span4Mux_v I__5390 (
            .O(N__23767),
            .I(N__23755));
    Span4Mux_h I__5389 (
            .O(N__23764),
            .I(N__23752));
    LocalMux I__5388 (
            .O(N__23761),
            .I(N__23749));
    LocalMux I__5387 (
            .O(N__23758),
            .I(N__23746));
    Span4Mux_h I__5386 (
            .O(N__23755),
            .I(N__23743));
    Span4Mux_h I__5385 (
            .O(N__23752),
            .I(N__23740));
    Span4Mux_v I__5384 (
            .O(N__23749),
            .I(N__23737));
    Span4Mux_h I__5383 (
            .O(N__23746),
            .I(N__23734));
    Odrv4 I__5382 (
            .O(N__23743),
            .I(\demux.N_417_i_0_o2Z0Z_9 ));
    Odrv4 I__5381 (
            .O(N__23740),
            .I(\demux.N_417_i_0_o2Z0Z_9 ));
    Odrv4 I__5380 (
            .O(N__23737),
            .I(\demux.N_417_i_0_o2Z0Z_9 ));
    Odrv4 I__5379 (
            .O(N__23734),
            .I(\demux.N_417_i_0_o2Z0Z_9 ));
    CascadeMux I__5378 (
            .O(N__23725),
            .I(N__23722));
    InMux I__5377 (
            .O(N__23722),
            .I(N__23718));
    InMux I__5376 (
            .O(N__23721),
            .I(N__23715));
    LocalMux I__5375 (
            .O(N__23718),
            .I(N__23709));
    LocalMux I__5374 (
            .O(N__23715),
            .I(N__23709));
    InMux I__5373 (
            .O(N__23714),
            .I(N__23706));
    Odrv4 I__5372 (
            .O(N__23709),
            .I(\demux.N_888 ));
    LocalMux I__5371 (
            .O(N__23706),
            .I(\demux.N_888 ));
    CascadeMux I__5370 (
            .O(N__23701),
            .I(N__23695));
    CascadeMux I__5369 (
            .O(N__23700),
            .I(N__23692));
    InMux I__5368 (
            .O(N__23699),
            .I(N__23689));
    InMux I__5367 (
            .O(N__23698),
            .I(N__23686));
    InMux I__5366 (
            .O(N__23695),
            .I(N__23683));
    InMux I__5365 (
            .O(N__23692),
            .I(N__23680));
    LocalMux I__5364 (
            .O(N__23689),
            .I(\demux.N_417_i_0_o2Z0Z_7 ));
    LocalMux I__5363 (
            .O(N__23686),
            .I(\demux.N_417_i_0_o2Z0Z_7 ));
    LocalMux I__5362 (
            .O(N__23683),
            .I(\demux.N_417_i_0_o2Z0Z_7 ));
    LocalMux I__5361 (
            .O(N__23680),
            .I(\demux.N_417_i_0_o2Z0Z_7 ));
    InMux I__5360 (
            .O(N__23671),
            .I(N__23668));
    LocalMux I__5359 (
            .O(N__23668),
            .I(N__23665));
    Span12Mux_s5_h I__5358 (
            .O(N__23665),
            .I(N__23662));
    Odrv12 I__5357 (
            .O(N__23662),
            .I(miso_data_in_7));
    InMux I__5356 (
            .O(N__23659),
            .I(N__23655));
    CascadeMux I__5355 (
            .O(N__23658),
            .I(N__23652));
    LocalMux I__5354 (
            .O(N__23655),
            .I(N__23649));
    InMux I__5353 (
            .O(N__23652),
            .I(N__23646));
    Span4Mux_v I__5352 (
            .O(N__23649),
            .I(N__23642));
    LocalMux I__5351 (
            .O(N__23646),
            .I(N__23639));
    InMux I__5350 (
            .O(N__23645),
            .I(N__23636));
    Odrv4 I__5349 (
            .O(N__23642),
            .I(\demux.N_874 ));
    Odrv12 I__5348 (
            .O(N__23639),
            .I(\demux.N_874 ));
    LocalMux I__5347 (
            .O(N__23636),
            .I(\demux.N_874 ));
    InMux I__5346 (
            .O(N__23629),
            .I(N__23626));
    LocalMux I__5345 (
            .O(N__23626),
            .I(N__23622));
    InMux I__5344 (
            .O(N__23625),
            .I(N__23619));
    Span4Mux_v I__5343 (
            .O(N__23622),
            .I(N__23612));
    LocalMux I__5342 (
            .O(N__23619),
            .I(N__23612));
    InMux I__5341 (
            .O(N__23618),
            .I(N__23609));
    InMux I__5340 (
            .O(N__23617),
            .I(N__23606));
    Odrv4 I__5339 (
            .O(N__23612),
            .I(\demux.N_418_i_0_o2Z0Z_8 ));
    LocalMux I__5338 (
            .O(N__23609),
            .I(\demux.N_418_i_0_o2Z0Z_8 ));
    LocalMux I__5337 (
            .O(N__23606),
            .I(\demux.N_418_i_0_o2Z0Z_8 ));
    CascadeMux I__5336 (
            .O(N__23599),
            .I(N__23596));
    InMux I__5335 (
            .O(N__23596),
            .I(N__23592));
    InMux I__5334 (
            .O(N__23595),
            .I(N__23589));
    LocalMux I__5333 (
            .O(N__23592),
            .I(N__23583));
    LocalMux I__5332 (
            .O(N__23589),
            .I(N__23583));
    CascadeMux I__5331 (
            .O(N__23588),
            .I(N__23579));
    Span4Mux_v I__5330 (
            .O(N__23583),
            .I(N__23576));
    InMux I__5329 (
            .O(N__23582),
            .I(N__23573));
    InMux I__5328 (
            .O(N__23579),
            .I(N__23570));
    Sp12to4 I__5327 (
            .O(N__23576),
            .I(N__23563));
    LocalMux I__5326 (
            .O(N__23573),
            .I(N__23563));
    LocalMux I__5325 (
            .O(N__23570),
            .I(N__23563));
    Odrv12 I__5324 (
            .O(N__23563),
            .I(\demux.N_418_i_0_o2Z0Z_9 ));
    InMux I__5323 (
            .O(N__23560),
            .I(N__23555));
    InMux I__5322 (
            .O(N__23559),
            .I(N__23552));
    InMux I__5321 (
            .O(N__23558),
            .I(N__23548));
    LocalMux I__5320 (
            .O(N__23555),
            .I(N__23543));
    LocalMux I__5319 (
            .O(N__23552),
            .I(N__23543));
    InMux I__5318 (
            .O(N__23551),
            .I(N__23540));
    LocalMux I__5317 (
            .O(N__23548),
            .I(\demux.N_418_i_0_o2Z0Z_7 ));
    Odrv4 I__5316 (
            .O(N__23543),
            .I(\demux.N_418_i_0_o2Z0Z_7 ));
    LocalMux I__5315 (
            .O(N__23540),
            .I(\demux.N_418_i_0_o2Z0Z_7 ));
    InMux I__5314 (
            .O(N__23533),
            .I(N__23530));
    LocalMux I__5313 (
            .O(N__23530),
            .I(N__23527));
    Odrv12 I__5312 (
            .O(N__23527),
            .I(miso_data_in_6));
    InMux I__5311 (
            .O(N__23524),
            .I(N__23521));
    LocalMux I__5310 (
            .O(N__23521),
            .I(N__23518));
    Span4Mux_h I__5309 (
            .O(N__23518),
            .I(N__23515));
    Odrv4 I__5308 (
            .O(N__23515),
            .I(demux_data_in_14));
    InMux I__5307 (
            .O(N__23512),
            .I(N__23509));
    LocalMux I__5306 (
            .O(N__23509),
            .I(\demux.N_880 ));
    InMux I__5305 (
            .O(N__23506),
            .I(N__23503));
    LocalMux I__5304 (
            .O(N__23503),
            .I(N__23500));
    Span4Mux_h I__5303 (
            .O(N__23500),
            .I(N__23497));
    Span4Mux_h I__5302 (
            .O(N__23497),
            .I(N__23494));
    Span4Mux_v I__5301 (
            .O(N__23494),
            .I(N__23491));
    Odrv4 I__5300 (
            .O(N__23491),
            .I(demux_data_in_36));
    InMux I__5299 (
            .O(N__23488),
            .I(N__23482));
    InMux I__5298 (
            .O(N__23487),
            .I(N__23482));
    LocalMux I__5297 (
            .O(N__23482),
            .I(N__23474));
    InMux I__5296 (
            .O(N__23481),
            .I(N__23469));
    InMux I__5295 (
            .O(N__23480),
            .I(N__23469));
    InMux I__5294 (
            .O(N__23479),
            .I(N__23466));
    InMux I__5293 (
            .O(N__23478),
            .I(N__23461));
    InMux I__5292 (
            .O(N__23477),
            .I(N__23461));
    Span4Mux_v I__5291 (
            .O(N__23474),
            .I(N__23456));
    LocalMux I__5290 (
            .O(N__23469),
            .I(N__23456));
    LocalMux I__5289 (
            .O(N__23466),
            .I(N__23453));
    LocalMux I__5288 (
            .O(N__23461),
            .I(N__23449));
    Span4Mux_h I__5287 (
            .O(N__23456),
            .I(N__23444));
    Span4Mux_h I__5286 (
            .O(N__23453),
            .I(N__23444));
    InMux I__5285 (
            .O(N__23452),
            .I(N__23441));
    Odrv4 I__5284 (
            .O(N__23449),
            .I(\demux.N_424_i_0_a2Z0Z_4 ));
    Odrv4 I__5283 (
            .O(N__23444),
            .I(\demux.N_424_i_0_a2Z0Z_4 ));
    LocalMux I__5282 (
            .O(N__23441),
            .I(\demux.N_424_i_0_a2Z0Z_4 ));
    CascadeMux I__5281 (
            .O(N__23434),
            .I(N__23430));
    CascadeMux I__5280 (
            .O(N__23433),
            .I(N__23427));
    InMux I__5279 (
            .O(N__23430),
            .I(N__23419));
    InMux I__5278 (
            .O(N__23427),
            .I(N__23419));
    CascadeMux I__5277 (
            .O(N__23426),
            .I(N__23416));
    CascadeMux I__5276 (
            .O(N__23425),
            .I(N__23413));
    CascadeMux I__5275 (
            .O(N__23424),
            .I(N__23409));
    LocalMux I__5274 (
            .O(N__23419),
            .I(N__23405));
    InMux I__5273 (
            .O(N__23416),
            .I(N__23400));
    InMux I__5272 (
            .O(N__23413),
            .I(N__23400));
    InMux I__5271 (
            .O(N__23412),
            .I(N__23397));
    InMux I__5270 (
            .O(N__23409),
            .I(N__23392));
    InMux I__5269 (
            .O(N__23408),
            .I(N__23392));
    Span4Mux_h I__5268 (
            .O(N__23405),
            .I(N__23387));
    LocalMux I__5267 (
            .O(N__23400),
            .I(N__23387));
    LocalMux I__5266 (
            .O(N__23397),
            .I(N__23384));
    LocalMux I__5265 (
            .O(N__23392),
            .I(\demux.N_424_i_0_a2Z0Z_5 ));
    Odrv4 I__5264 (
            .O(N__23387),
            .I(\demux.N_424_i_0_a2Z0Z_5 ));
    Odrv4 I__5263 (
            .O(N__23384),
            .I(\demux.N_424_i_0_a2Z0Z_5 ));
    InMux I__5262 (
            .O(N__23377),
            .I(N__23374));
    LocalMux I__5261 (
            .O(N__23374),
            .I(demux_data_in_108));
    InMux I__5260 (
            .O(N__23371),
            .I(N__23362));
    InMux I__5259 (
            .O(N__23370),
            .I(N__23357));
    InMux I__5258 (
            .O(N__23369),
            .I(N__23357));
    InMux I__5257 (
            .O(N__23368),
            .I(N__23352));
    InMux I__5256 (
            .O(N__23367),
            .I(N__23352));
    InMux I__5255 (
            .O(N__23366),
            .I(N__23347));
    InMux I__5254 (
            .O(N__23365),
            .I(N__23347));
    LocalMux I__5253 (
            .O(N__23362),
            .I(N__23343));
    LocalMux I__5252 (
            .O(N__23357),
            .I(N__23340));
    LocalMux I__5251 (
            .O(N__23352),
            .I(N__23335));
    LocalMux I__5250 (
            .O(N__23347),
            .I(N__23335));
    InMux I__5249 (
            .O(N__23346),
            .I(N__23332));
    Span4Mux_h I__5248 (
            .O(N__23343),
            .I(N__23327));
    Span4Mux_h I__5247 (
            .O(N__23340),
            .I(N__23327));
    Span4Mux_h I__5246 (
            .O(N__23335),
            .I(N__23324));
    LocalMux I__5245 (
            .O(N__23332),
            .I(\demux.N_424_i_0_a2Z0Z_11 ));
    Odrv4 I__5244 (
            .O(N__23327),
            .I(\demux.N_424_i_0_a2Z0Z_11 ));
    Odrv4 I__5243 (
            .O(N__23324),
            .I(\demux.N_424_i_0_a2Z0Z_11 ));
    CascadeMux I__5242 (
            .O(N__23317),
            .I(\demux.N_420_i_0_o2Z0Z_0_cascade_ ));
    InMux I__5241 (
            .O(N__23314),
            .I(N__23311));
    LocalMux I__5240 (
            .O(N__23311),
            .I(N__23308));
    Span4Mux_h I__5239 (
            .O(N__23308),
            .I(N__23305));
    Odrv4 I__5238 (
            .O(N__23305),
            .I(demux_data_in_92));
    InMux I__5237 (
            .O(N__23302),
            .I(N__23299));
    LocalMux I__5236 (
            .O(N__23299),
            .I(N__23290));
    InMux I__5235 (
            .O(N__23298),
            .I(N__23287));
    InMux I__5234 (
            .O(N__23297),
            .I(N__23284));
    InMux I__5233 (
            .O(N__23296),
            .I(N__23281));
    InMux I__5232 (
            .O(N__23295),
            .I(N__23278));
    InMux I__5231 (
            .O(N__23294),
            .I(N__23273));
    InMux I__5230 (
            .O(N__23293),
            .I(N__23273));
    Span4Mux_h I__5229 (
            .O(N__23290),
            .I(N__23267));
    LocalMux I__5228 (
            .O(N__23287),
            .I(N__23267));
    LocalMux I__5227 (
            .O(N__23284),
            .I(N__23264));
    LocalMux I__5226 (
            .O(N__23281),
            .I(N__23257));
    LocalMux I__5225 (
            .O(N__23278),
            .I(N__23257));
    LocalMux I__5224 (
            .O(N__23273),
            .I(N__23257));
    InMux I__5223 (
            .O(N__23272),
            .I(N__23254));
    Span4Mux_v I__5222 (
            .O(N__23267),
            .I(N__23251));
    Span4Mux_h I__5221 (
            .O(N__23264),
            .I(N__23248));
    Span4Mux_v I__5220 (
            .O(N__23257),
            .I(N__23243));
    LocalMux I__5219 (
            .O(N__23254),
            .I(N__23243));
    Odrv4 I__5218 (
            .O(N__23251),
            .I(\demux.N_424_i_0_a2Z0Z_2 ));
    Odrv4 I__5217 (
            .O(N__23248),
            .I(\demux.N_424_i_0_a2Z0Z_2 ));
    Odrv4 I__5216 (
            .O(N__23243),
            .I(\demux.N_424_i_0_a2Z0Z_2 ));
    InMux I__5215 (
            .O(N__23236),
            .I(N__23233));
    LocalMux I__5214 (
            .O(N__23233),
            .I(N__23230));
    Span4Mux_v I__5213 (
            .O(N__23230),
            .I(N__23227));
    Span4Mux_s3_h I__5212 (
            .O(N__23227),
            .I(N__23224));
    Odrv4 I__5211 (
            .O(N__23224),
            .I(demux_data_in_12));
    CascadeMux I__5210 (
            .O(N__23221),
            .I(\demux.N_420_i_0_o2Z0Z_1_cascade_ ));
    InMux I__5209 (
            .O(N__23218),
            .I(N__23215));
    LocalMux I__5208 (
            .O(N__23215),
            .I(N__23212));
    Odrv4 I__5207 (
            .O(N__23212),
            .I(\demux.N_420_i_0_a3Z0Z_4 ));
    InMux I__5206 (
            .O(N__23209),
            .I(N__23206));
    LocalMux I__5205 (
            .O(N__23206),
            .I(N__23203));
    Sp12to4 I__5204 (
            .O(N__23203),
            .I(N__23200));
    Odrv12 I__5203 (
            .O(N__23200),
            .I(demux_data_in_7));
    CascadeMux I__5202 (
            .O(N__23197),
            .I(\demux.N_888_cascade_ ));
    InMux I__5201 (
            .O(N__23194),
            .I(N__23191));
    LocalMux I__5200 (
            .O(N__23191),
            .I(N__23188));
    Sp12to4 I__5199 (
            .O(N__23188),
            .I(N__23185));
    Odrv12 I__5198 (
            .O(N__23185),
            .I(demux_data_in_6));
    InMux I__5197 (
            .O(N__23182),
            .I(N__23179));
    LocalMux I__5196 (
            .O(N__23179),
            .I(N__23176));
    Odrv4 I__5195 (
            .O(N__23176),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_0 ));
    InMux I__5194 (
            .O(N__23173),
            .I(N__23170));
    LocalMux I__5193 (
            .O(N__23170),
            .I(N__23167));
    Odrv4 I__5192 (
            .O(N__23167),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_10 ));
    InMux I__5191 (
            .O(N__23164),
            .I(N__23161));
    LocalMux I__5190 (
            .O(N__23161),
            .I(N__23158));
    Odrv4 I__5189 (
            .O(N__23158),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_12 ));
    InMux I__5188 (
            .O(N__23155),
            .I(N__23152));
    LocalMux I__5187 (
            .O(N__23152),
            .I(N__23149));
    Odrv4 I__5186 (
            .O(N__23149),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_18 ));
    InMux I__5185 (
            .O(N__23146),
            .I(N__23143));
    LocalMux I__5184 (
            .O(N__23143),
            .I(N__23140));
    Span4Mux_h I__5183 (
            .O(N__23140),
            .I(N__23137));
    Odrv4 I__5182 (
            .O(N__23137),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_15 ));
    InMux I__5181 (
            .O(N__23134),
            .I(N__23131));
    LocalMux I__5180 (
            .O(N__23131),
            .I(N__23128));
    Odrv4 I__5179 (
            .O(N__23128),
            .I(\sb_translator_1.rgb_data_tmpZ0Z_16 ));
    InMux I__5178 (
            .O(N__23125),
            .I(N__23122));
    LocalMux I__5177 (
            .O(N__23122),
            .I(N__23119));
    Odrv4 I__5176 (
            .O(N__23119),
            .I(demux_data_in_94));
    InMux I__5175 (
            .O(N__23116),
            .I(N__23113));
    LocalMux I__5174 (
            .O(N__23113),
            .I(demux_data_in_110));
    CascadeMux I__5173 (
            .O(N__23110),
            .I(\demux.N_418_i_0_o2Z0Z_0_cascade_ ));
    InMux I__5172 (
            .O(N__23107),
            .I(N__23104));
    LocalMux I__5171 (
            .O(N__23104),
            .I(N__23101));
    Span4Mux_h I__5170 (
            .O(N__23101),
            .I(N__23098));
    Span4Mux_h I__5169 (
            .O(N__23098),
            .I(N__23095));
    Span4Mux_v I__5168 (
            .O(N__23095),
            .I(N__23092));
    Odrv4 I__5167 (
            .O(N__23092),
            .I(demux_data_in_38));
    InMux I__5166 (
            .O(N__23089),
            .I(N__23086));
    LocalMux I__5165 (
            .O(N__23086),
            .I(N__23083));
    Span12Mux_s10_h I__5164 (
            .O(N__23083),
            .I(N__23080));
    Odrv12 I__5163 (
            .O(N__23080),
            .I(demux_data_in_46));
    CascadeMux I__5162 (
            .O(N__23077),
            .I(\demux.N_418_i_0_o2Z0Z_1_cascade_ ));
    InMux I__5161 (
            .O(N__23074),
            .I(N__23068));
    InMux I__5160 (
            .O(N__23073),
            .I(N__23065));
    InMux I__5159 (
            .O(N__23072),
            .I(N__23061));
    InMux I__5158 (
            .O(N__23071),
            .I(N__23058));
    LocalMux I__5157 (
            .O(N__23068),
            .I(N__23050));
    LocalMux I__5156 (
            .O(N__23065),
            .I(N__23050));
    InMux I__5155 (
            .O(N__23064),
            .I(N__23047));
    LocalMux I__5154 (
            .O(N__23061),
            .I(N__23042));
    LocalMux I__5153 (
            .O(N__23058),
            .I(N__23042));
    InMux I__5152 (
            .O(N__23057),
            .I(N__23037));
    InMux I__5151 (
            .O(N__23056),
            .I(N__23037));
    InMux I__5150 (
            .O(N__23055),
            .I(N__23034));
    Span4Mux_h I__5149 (
            .O(N__23050),
            .I(N__23031));
    LocalMux I__5148 (
            .O(N__23047),
            .I(N__23028));
    Span4Mux_v I__5147 (
            .O(N__23042),
            .I(N__23023));
    LocalMux I__5146 (
            .O(N__23037),
            .I(N__23023));
    LocalMux I__5145 (
            .O(N__23034),
            .I(N__23020));
    Odrv4 I__5144 (
            .O(N__23031),
            .I(\demux.N_424_i_0_a2Z0Z_8 ));
    Odrv4 I__5143 (
            .O(N__23028),
            .I(\demux.N_424_i_0_a2Z0Z_8 ));
    Odrv4 I__5142 (
            .O(N__23023),
            .I(\demux.N_424_i_0_a2Z0Z_8 ));
    Odrv4 I__5141 (
            .O(N__23020),
            .I(\demux.N_424_i_0_a2Z0Z_8 ));
    InMux I__5140 (
            .O(N__23011),
            .I(N__23005));
    InMux I__5139 (
            .O(N__23010),
            .I(N__23000));
    InMux I__5138 (
            .O(N__23009),
            .I(N__23000));
    InMux I__5137 (
            .O(N__23008),
            .I(N__22994));
    LocalMux I__5136 (
            .O(N__23005),
            .I(N__22991));
    LocalMux I__5135 (
            .O(N__23000),
            .I(N__22988));
    InMux I__5134 (
            .O(N__22999),
            .I(N__22981));
    InMux I__5133 (
            .O(N__22998),
            .I(N__22981));
    InMux I__5132 (
            .O(N__22997),
            .I(N__22981));
    LocalMux I__5131 (
            .O(N__22994),
            .I(N__22975));
    Span4Mux_h I__5130 (
            .O(N__22991),
            .I(N__22972));
    Span4Mux_h I__5129 (
            .O(N__22988),
            .I(N__22969));
    LocalMux I__5128 (
            .O(N__22981),
            .I(N__22966));
    InMux I__5127 (
            .O(N__22980),
            .I(N__22959));
    InMux I__5126 (
            .O(N__22979),
            .I(N__22959));
    InMux I__5125 (
            .O(N__22978),
            .I(N__22959));
    Span4Mux_v I__5124 (
            .O(N__22975),
            .I(N__22954));
    Span4Mux_h I__5123 (
            .O(N__22972),
            .I(N__22954));
    Odrv4 I__5122 (
            .O(N__22969),
            .I(\sb_translator_1.stateZ0Z_6 ));
    Odrv12 I__5121 (
            .O(N__22966),
            .I(\sb_translator_1.stateZ0Z_6 ));
    LocalMux I__5120 (
            .O(N__22959),
            .I(\sb_translator_1.stateZ0Z_6 ));
    Odrv4 I__5119 (
            .O(N__22954),
            .I(\sb_translator_1.stateZ0Z_6 ));
    InMux I__5118 (
            .O(N__22945),
            .I(N__22941));
    InMux I__5117 (
            .O(N__22944),
            .I(N__22938));
    LocalMux I__5116 (
            .O(N__22941),
            .I(N__22933));
    LocalMux I__5115 (
            .O(N__22938),
            .I(N__22933));
    Span4Mux_v I__5114 (
            .O(N__22933),
            .I(N__22930));
    Odrv4 I__5113 (
            .O(N__22930),
            .I(mosi_data_out_15));
    InMux I__5112 (
            .O(N__22927),
            .I(N__22923));
    InMux I__5111 (
            .O(N__22926),
            .I(N__22920));
    LocalMux I__5110 (
            .O(N__22923),
            .I(N__22916));
    LocalMux I__5109 (
            .O(N__22920),
            .I(N__22913));
    InMux I__5108 (
            .O(N__22919),
            .I(N__22910));
    Span4Mux_s2_h I__5107 (
            .O(N__22916),
            .I(N__22907));
    Odrv12 I__5106 (
            .O(N__22913),
            .I(\sb_translator_1.cntZ0Z_7 ));
    LocalMux I__5105 (
            .O(N__22910),
            .I(\sb_translator_1.cntZ0Z_7 ));
    Odrv4 I__5104 (
            .O(N__22907),
            .I(\sb_translator_1.cntZ0Z_7 ));
    CascadeMux I__5103 (
            .O(N__22900),
            .I(N__22897));
    InMux I__5102 (
            .O(N__22897),
            .I(N__22894));
    LocalMux I__5101 (
            .O(N__22894),
            .I(N__22891));
    Odrv4 I__5100 (
            .O(N__22891),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_7 ));
    InMux I__5099 (
            .O(N__22888),
            .I(N__22885));
    LocalMux I__5098 (
            .O(N__22885),
            .I(N__22882));
    Span4Mux_v I__5097 (
            .O(N__22882),
            .I(N__22879));
    Odrv4 I__5096 (
            .O(N__22879),
            .I(\ws2812.new_data_req_e_1 ));
    CascadeMux I__5095 (
            .O(N__22876),
            .I(\ws2812.N_140_cascade_ ));
    InMux I__5094 (
            .O(N__22873),
            .I(N__22870));
    LocalMux I__5093 (
            .O(N__22870),
            .I(N__22866));
    InMux I__5092 (
            .O(N__22869),
            .I(N__22863));
    Span12Mux_s8_v I__5091 (
            .O(N__22866),
            .I(N__22860));
    LocalMux I__5090 (
            .O(N__22863),
            .I(ws2812_next_led));
    Odrv12 I__5089 (
            .O(N__22860),
            .I(ws2812_next_led));
    InMux I__5088 (
            .O(N__22855),
            .I(N__22852));
    LocalMux I__5087 (
            .O(N__22852),
            .I(\sb_translator_1.state56_a_5_8 ));
    InMux I__5086 (
            .O(N__22849),
            .I(N__22846));
    LocalMux I__5085 (
            .O(N__22846),
            .I(\sb_translator_1.state56_a_5_9 ));
    CascadeMux I__5084 (
            .O(N__22843),
            .I(\sb_translator_1.N_318_i_i_o2_11_cascade_ ));
    InMux I__5083 (
            .O(N__22840),
            .I(N__22837));
    LocalMux I__5082 (
            .O(N__22837),
            .I(\sb_translator_1.state56_a_5_15 ));
    InMux I__5081 (
            .O(N__22834),
            .I(N__22831));
    LocalMux I__5080 (
            .O(N__22831),
            .I(\sb_translator_1.N_318_i_i_o2_14 ));
    CascadeMux I__5079 (
            .O(N__22828),
            .I(N__22825));
    InMux I__5078 (
            .O(N__22825),
            .I(N__22822));
    LocalMux I__5077 (
            .O(N__22822),
            .I(N__22817));
    InMux I__5076 (
            .O(N__22821),
            .I(N__22812));
    InMux I__5075 (
            .O(N__22820),
            .I(N__22812));
    Span4Mux_s3_v I__5074 (
            .O(N__22817),
            .I(N__22807));
    LocalMux I__5073 (
            .O(N__22812),
            .I(N__22807));
    Span4Mux_h I__5072 (
            .O(N__22807),
            .I(N__22804));
    Span4Mux_v I__5071 (
            .O(N__22804),
            .I(N__22801));
    Odrv4 I__5070 (
            .O(N__22801),
            .I(\sb_translator_1.state_RNII30CZ0Z_0 ));
    IoInMux I__5069 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__5068 (
            .O(N__22795),
            .I(N__22792));
    Odrv4 I__5067 (
            .O(N__22792),
            .I(\sb_translator_1.stateZ0Z_1 ));
    CascadeMux I__5066 (
            .O(N__22789),
            .I(N__22776));
    CascadeMux I__5065 (
            .O(N__22788),
            .I(N__22773));
    CascadeMux I__5064 (
            .O(N__22787),
            .I(N__22770));
    CascadeMux I__5063 (
            .O(N__22786),
            .I(N__22767));
    InMux I__5062 (
            .O(N__22785),
            .I(N__22756));
    CascadeMux I__5061 (
            .O(N__22784),
            .I(N__22753));
    CascadeMux I__5060 (
            .O(N__22783),
            .I(N__22748));
    CascadeMux I__5059 (
            .O(N__22782),
            .I(N__22745));
    CascadeMux I__5058 (
            .O(N__22781),
            .I(N__22742));
    CascadeMux I__5057 (
            .O(N__22780),
            .I(N__22739));
    CascadeMux I__5056 (
            .O(N__22779),
            .I(N__22736));
    InMux I__5055 (
            .O(N__22776),
            .I(N__22725));
    InMux I__5054 (
            .O(N__22773),
            .I(N__22725));
    InMux I__5053 (
            .O(N__22770),
            .I(N__22725));
    InMux I__5052 (
            .O(N__22767),
            .I(N__22725));
    InMux I__5051 (
            .O(N__22766),
            .I(N__22716));
    InMux I__5050 (
            .O(N__22765),
            .I(N__22716));
    InMux I__5049 (
            .O(N__22764),
            .I(N__22716));
    InMux I__5048 (
            .O(N__22763),
            .I(N__22716));
    InMux I__5047 (
            .O(N__22762),
            .I(N__22713));
    InMux I__5046 (
            .O(N__22761),
            .I(N__22706));
    InMux I__5045 (
            .O(N__22760),
            .I(N__22706));
    InMux I__5044 (
            .O(N__22759),
            .I(N__22706));
    LocalMux I__5043 (
            .O(N__22756),
            .I(N__22703));
    InMux I__5042 (
            .O(N__22753),
            .I(N__22696));
    InMux I__5041 (
            .O(N__22752),
            .I(N__22696));
    InMux I__5040 (
            .O(N__22751),
            .I(N__22696));
    InMux I__5039 (
            .O(N__22748),
            .I(N__22691));
    InMux I__5038 (
            .O(N__22745),
            .I(N__22691));
    InMux I__5037 (
            .O(N__22742),
            .I(N__22680));
    InMux I__5036 (
            .O(N__22739),
            .I(N__22680));
    InMux I__5035 (
            .O(N__22736),
            .I(N__22680));
    InMux I__5034 (
            .O(N__22735),
            .I(N__22680));
    InMux I__5033 (
            .O(N__22734),
            .I(N__22680));
    LocalMux I__5032 (
            .O(N__22725),
            .I(N__22671));
    LocalMux I__5031 (
            .O(N__22716),
            .I(N__22671));
    LocalMux I__5030 (
            .O(N__22713),
            .I(N__22671));
    LocalMux I__5029 (
            .O(N__22706),
            .I(N__22671));
    Span4Mux_v I__5028 (
            .O(N__22703),
            .I(N__22668));
    LocalMux I__5027 (
            .O(N__22696),
            .I(N__22665));
    LocalMux I__5026 (
            .O(N__22691),
            .I(N__22662));
    LocalMux I__5025 (
            .O(N__22680),
            .I(N__22659));
    Span4Mux_v I__5024 (
            .O(N__22671),
            .I(N__22652));
    Span4Mux_v I__5023 (
            .O(N__22668),
            .I(N__22652));
    Span4Mux_h I__5022 (
            .O(N__22665),
            .I(N__22652));
    Odrv12 I__5021 (
            .O(N__22662),
            .I(mosi_data_out_23));
    Odrv4 I__5020 (
            .O(N__22659),
            .I(mosi_data_out_23));
    Odrv4 I__5019 (
            .O(N__22652),
            .I(mosi_data_out_23));
    CascadeMux I__5018 (
            .O(N__22645),
            .I(N__22640));
    InMux I__5017 (
            .O(N__22644),
            .I(N__22635));
    InMux I__5016 (
            .O(N__22643),
            .I(N__22632));
    InMux I__5015 (
            .O(N__22640),
            .I(N__22629));
    InMux I__5014 (
            .O(N__22639),
            .I(N__22624));
    InMux I__5013 (
            .O(N__22638),
            .I(N__22624));
    LocalMux I__5012 (
            .O(N__22635),
            .I(N__22619));
    LocalMux I__5011 (
            .O(N__22632),
            .I(N__22619));
    LocalMux I__5010 (
            .O(N__22629),
            .I(N__22614));
    LocalMux I__5009 (
            .O(N__22624),
            .I(N__22614));
    Span4Mux_v I__5008 (
            .O(N__22619),
            .I(N__22611));
    Span12Mux_s9_h I__5007 (
            .O(N__22614),
            .I(N__22608));
    Odrv4 I__5006 (
            .O(N__22611),
            .I(mosi_data_out_21));
    Odrv12 I__5005 (
            .O(N__22608),
            .I(mosi_data_out_21));
    CascadeMux I__5004 (
            .O(N__22603),
            .I(N__22599));
    InMux I__5003 (
            .O(N__22602),
            .I(N__22591));
    InMux I__5002 (
            .O(N__22599),
            .I(N__22591));
    InMux I__5001 (
            .O(N__22598),
            .I(N__22591));
    LocalMux I__5000 (
            .O(N__22591),
            .I(N__22588));
    Span12Mux_s9_h I__4999 (
            .O(N__22588),
            .I(N__22585));
    Odrv12 I__4998 (
            .O(N__22585),
            .I(\sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0 ));
    InMux I__4997 (
            .O(N__22582),
            .I(N__22579));
    LocalMux I__4996 (
            .O(N__22579),
            .I(N__22575));
    InMux I__4995 (
            .O(N__22578),
            .I(N__22572));
    Span4Mux_h I__4994 (
            .O(N__22575),
            .I(N__22569));
    LocalMux I__4993 (
            .O(N__22572),
            .I(mosi_data_out_12));
    Odrv4 I__4992 (
            .O(N__22569),
            .I(mosi_data_out_12));
    InMux I__4991 (
            .O(N__22564),
            .I(N__22561));
    LocalMux I__4990 (
            .O(N__22561),
            .I(N__22557));
    InMux I__4989 (
            .O(N__22560),
            .I(N__22553));
    Span4Mux_h I__4988 (
            .O(N__22557),
            .I(N__22550));
    InMux I__4987 (
            .O(N__22556),
            .I(N__22547));
    LocalMux I__4986 (
            .O(N__22553),
            .I(N__22544));
    Odrv4 I__4985 (
            .O(N__22550),
            .I(\sb_translator_1.cntZ0Z_4 ));
    LocalMux I__4984 (
            .O(N__22547),
            .I(\sb_translator_1.cntZ0Z_4 ));
    Odrv4 I__4983 (
            .O(N__22544),
            .I(\sb_translator_1.cntZ0Z_4 ));
    InMux I__4982 (
            .O(N__22537),
            .I(N__22534));
    LocalMux I__4981 (
            .O(N__22534),
            .I(N__22531));
    Span4Mux_h I__4980 (
            .O(N__22531),
            .I(N__22528));
    Odrv4 I__4979 (
            .O(N__22528),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_4 ));
    InMux I__4978 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__4977 (
            .O(N__22522),
            .I(N__22518));
    InMux I__4976 (
            .O(N__22521),
            .I(N__22515));
    Span4Mux_h I__4975 (
            .O(N__22518),
            .I(N__22512));
    LocalMux I__4974 (
            .O(N__22515),
            .I(mosi_data_out_14));
    Odrv4 I__4973 (
            .O(N__22512),
            .I(mosi_data_out_14));
    InMux I__4972 (
            .O(N__22507),
            .I(N__22503));
    InMux I__4971 (
            .O(N__22506),
            .I(N__22499));
    LocalMux I__4970 (
            .O(N__22503),
            .I(N__22496));
    InMux I__4969 (
            .O(N__22502),
            .I(N__22493));
    LocalMux I__4968 (
            .O(N__22499),
            .I(N__22490));
    Odrv12 I__4967 (
            .O(N__22496),
            .I(\sb_translator_1.cntZ0Z_6 ));
    LocalMux I__4966 (
            .O(N__22493),
            .I(\sb_translator_1.cntZ0Z_6 ));
    Odrv4 I__4965 (
            .O(N__22490),
            .I(\sb_translator_1.cntZ0Z_6 ));
    InMux I__4964 (
            .O(N__22483),
            .I(N__22480));
    LocalMux I__4963 (
            .O(N__22480),
            .I(N__22477));
    Span4Mux_h I__4962 (
            .O(N__22477),
            .I(N__22474));
    Odrv4 I__4961 (
            .O(N__22474),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_6 ));
    InMux I__4960 (
            .O(N__22471),
            .I(N__22468));
    LocalMux I__4959 (
            .O(N__22468),
            .I(\sb_translator_1.state56_a_5_6 ));
    InMux I__4958 (
            .O(N__22465),
            .I(N__22462));
    LocalMux I__4957 (
            .O(N__22462),
            .I(\sb_translator_1.state56_a_5_11 ));
    CascadeMux I__4956 (
            .O(N__22459),
            .I(N__22456));
    InMux I__4955 (
            .O(N__22456),
            .I(N__22453));
    LocalMux I__4954 (
            .O(N__22453),
            .I(\sb_translator_1.state56_a_5_5 ));
    InMux I__4953 (
            .O(N__22450),
            .I(N__22447));
    LocalMux I__4952 (
            .O(N__22447),
            .I(\sb_translator_1.state56_a_5_13 ));
    InMux I__4951 (
            .O(N__22444),
            .I(N__22441));
    LocalMux I__4950 (
            .O(N__22441),
            .I(\sb_translator_1.state56_a_5_14 ));
    CascadeMux I__4949 (
            .O(N__22438),
            .I(\sb_translator_1.N_318_i_i_o2_12_cascade_ ));
    InMux I__4948 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__4947 (
            .O(N__22432),
            .I(N__22429));
    Odrv4 I__4946 (
            .O(N__22429),
            .I(\sb_translator_1.state56_17 ));
    InMux I__4945 (
            .O(N__22426),
            .I(N__22423));
    LocalMux I__4944 (
            .O(N__22423),
            .I(N__22418));
    InMux I__4943 (
            .O(N__22422),
            .I(N__22412));
    InMux I__4942 (
            .O(N__22421),
            .I(N__22412));
    Span4Mux_s3_v I__4941 (
            .O(N__22418),
            .I(N__22409));
    InMux I__4940 (
            .O(N__22417),
            .I(N__22406));
    LocalMux I__4939 (
            .O(N__22412),
            .I(N__22396));
    Span4Mux_v I__4938 (
            .O(N__22409),
            .I(N__22396));
    LocalMux I__4937 (
            .O(N__22406),
            .I(N__22393));
    InMux I__4936 (
            .O(N__22405),
            .I(N__22382));
    InMux I__4935 (
            .O(N__22404),
            .I(N__22382));
    InMux I__4934 (
            .O(N__22403),
            .I(N__22382));
    InMux I__4933 (
            .O(N__22402),
            .I(N__22382));
    InMux I__4932 (
            .O(N__22401),
            .I(N__22382));
    Span4Mux_h I__4931 (
            .O(N__22396),
            .I(N__22377));
    Span4Mux_h I__4930 (
            .O(N__22393),
            .I(N__22377));
    LocalMux I__4929 (
            .O(N__22382),
            .I(N__22374));
    Odrv4 I__4928 (
            .O(N__22377),
            .I(\sb_translator_1.state_leds_RNIGMAHZ0 ));
    Odrv12 I__4927 (
            .O(N__22374),
            .I(\sb_translator_1.state_leds_RNIGMAHZ0 ));
    CascadeMux I__4926 (
            .O(N__22369),
            .I(\sb_translator_1.N_318_i_i_o2_15_cascade_ ));
    CascadeMux I__4925 (
            .O(N__22366),
            .I(\sb_translator_1.N_712_cascade_ ));
    CEMux I__4924 (
            .O(N__22363),
            .I(N__22359));
    CEMux I__4923 (
            .O(N__22362),
            .I(N__22356));
    LocalMux I__4922 (
            .O(N__22359),
            .I(N__22350));
    LocalMux I__4921 (
            .O(N__22356),
            .I(N__22350));
    CEMux I__4920 (
            .O(N__22355),
            .I(N__22344));
    Span4Mux_v I__4919 (
            .O(N__22350),
            .I(N__22341));
    CEMux I__4918 (
            .O(N__22349),
            .I(N__22338));
    CEMux I__4917 (
            .O(N__22348),
            .I(N__22327));
    InMux I__4916 (
            .O(N__22347),
            .I(N__22315));
    LocalMux I__4915 (
            .O(N__22344),
            .I(N__22312));
    Span4Mux_s0_v I__4914 (
            .O(N__22341),
            .I(N__22307));
    LocalMux I__4913 (
            .O(N__22338),
            .I(N__22307));
    InMux I__4912 (
            .O(N__22337),
            .I(N__22296));
    InMux I__4911 (
            .O(N__22336),
            .I(N__22296));
    InMux I__4910 (
            .O(N__22335),
            .I(N__22296));
    InMux I__4909 (
            .O(N__22334),
            .I(N__22296));
    InMux I__4908 (
            .O(N__22333),
            .I(N__22287));
    InMux I__4907 (
            .O(N__22332),
            .I(N__22287));
    InMux I__4906 (
            .O(N__22331),
            .I(N__22287));
    InMux I__4905 (
            .O(N__22330),
            .I(N__22287));
    LocalMux I__4904 (
            .O(N__22327),
            .I(N__22284));
    InMux I__4903 (
            .O(N__22326),
            .I(N__22275));
    InMux I__4902 (
            .O(N__22325),
            .I(N__22275));
    InMux I__4901 (
            .O(N__22324),
            .I(N__22275));
    InMux I__4900 (
            .O(N__22323),
            .I(N__22275));
    InMux I__4899 (
            .O(N__22322),
            .I(N__22272));
    InMux I__4898 (
            .O(N__22321),
            .I(N__22263));
    InMux I__4897 (
            .O(N__22320),
            .I(N__22263));
    InMux I__4896 (
            .O(N__22319),
            .I(N__22263));
    InMux I__4895 (
            .O(N__22318),
            .I(N__22263));
    LocalMux I__4894 (
            .O(N__22315),
            .I(N__22260));
    Span4Mux_h I__4893 (
            .O(N__22312),
            .I(N__22254));
    Span4Mux_v I__4892 (
            .O(N__22307),
            .I(N__22254));
    InMux I__4891 (
            .O(N__22306),
            .I(N__22249));
    InMux I__4890 (
            .O(N__22305),
            .I(N__22249));
    LocalMux I__4889 (
            .O(N__22296),
            .I(N__22244));
    LocalMux I__4888 (
            .O(N__22287),
            .I(N__22244));
    Span4Mux_s2_v I__4887 (
            .O(N__22284),
            .I(N__22233));
    LocalMux I__4886 (
            .O(N__22275),
            .I(N__22233));
    LocalMux I__4885 (
            .O(N__22272),
            .I(N__22233));
    LocalMux I__4884 (
            .O(N__22263),
            .I(N__22233));
    Span4Mux_h I__4883 (
            .O(N__22260),
            .I(N__22233));
    InMux I__4882 (
            .O(N__22259),
            .I(N__22230));
    Span4Mux_v I__4881 (
            .O(N__22254),
            .I(N__22227));
    LocalMux I__4880 (
            .O(N__22249),
            .I(N__22220));
    Span4Mux_v I__4879 (
            .O(N__22244),
            .I(N__22220));
    Span4Mux_v I__4878 (
            .O(N__22233),
            .I(N__22220));
    LocalMux I__4877 (
            .O(N__22230),
            .I(N__22217));
    Odrv4 I__4876 (
            .O(N__22227),
            .I(\sb_translator_1.num_leds_1_sqmuxa ));
    Odrv4 I__4875 (
            .O(N__22220),
            .I(\sb_translator_1.num_leds_1_sqmuxa ));
    Odrv12 I__4874 (
            .O(N__22217),
            .I(\sb_translator_1.num_leds_1_sqmuxa ));
    CascadeMux I__4873 (
            .O(N__22210),
            .I(N__22207));
    InMux I__4872 (
            .O(N__22207),
            .I(N__22193));
    InMux I__4871 (
            .O(N__22206),
            .I(N__22176));
    InMux I__4870 (
            .O(N__22205),
            .I(N__22176));
    InMux I__4869 (
            .O(N__22204),
            .I(N__22176));
    InMux I__4868 (
            .O(N__22203),
            .I(N__22176));
    InMux I__4867 (
            .O(N__22202),
            .I(N__22176));
    InMux I__4866 (
            .O(N__22201),
            .I(N__22176));
    InMux I__4865 (
            .O(N__22200),
            .I(N__22176));
    InMux I__4864 (
            .O(N__22199),
            .I(N__22176));
    InMux I__4863 (
            .O(N__22198),
            .I(N__22169));
    InMux I__4862 (
            .O(N__22197),
            .I(N__22169));
    InMux I__4861 (
            .O(N__22196),
            .I(N__22169));
    LocalMux I__4860 (
            .O(N__22193),
            .I(N__22166));
    LocalMux I__4859 (
            .O(N__22176),
            .I(N__22163));
    LocalMux I__4858 (
            .O(N__22169),
            .I(N__22160));
    Span4Mux_v I__4857 (
            .O(N__22166),
            .I(N__22157));
    Span4Mux_v I__4856 (
            .O(N__22163),
            .I(N__22152));
    Span4Mux_v I__4855 (
            .O(N__22160),
            .I(N__22152));
    Span4Mux_h I__4854 (
            .O(N__22157),
            .I(N__22146));
    Span4Mux_v I__4853 (
            .O(N__22152),
            .I(N__22146));
    InMux I__4852 (
            .O(N__22151),
            .I(N__22143));
    Span4Mux_h I__4851 (
            .O(N__22146),
            .I(N__22140));
    LocalMux I__4850 (
            .O(N__22143),
            .I(\sb_translator_1.stateZ0Z_7 ));
    Odrv4 I__4849 (
            .O(N__22140),
            .I(\sb_translator_1.stateZ0Z_7 ));
    InMux I__4848 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__4847 (
            .O(N__22132),
            .I(\sb_translator_1.state56_a_5_2 ));
    InMux I__4846 (
            .O(N__22129),
            .I(N__22126));
    LocalMux I__4845 (
            .O(N__22126),
            .I(\sb_translator_1.state56_a_5_7 ));
    CascadeMux I__4844 (
            .O(N__22123),
            .I(N__22120));
    InMux I__4843 (
            .O(N__22120),
            .I(N__22117));
    LocalMux I__4842 (
            .O(N__22117),
            .I(N__22114));
    Odrv4 I__4841 (
            .O(N__22114),
            .I(\sb_translator_1.N_318_i_i_o2_0 ));
    InMux I__4840 (
            .O(N__22111),
            .I(N__22108));
    LocalMux I__4839 (
            .O(N__22108),
            .I(\sb_translator_1.state56_a_5_12 ));
    InMux I__4838 (
            .O(N__22105),
            .I(N__22102));
    LocalMux I__4837 (
            .O(N__22102),
            .I(\sb_translator_1.N_318_i_i_o2_8 ));
    InMux I__4836 (
            .O(N__22099),
            .I(N__22096));
    LocalMux I__4835 (
            .O(N__22096),
            .I(N__22093));
    Span4Mux_s3_v I__4834 (
            .O(N__22093),
            .I(N__22090));
    Span4Mux_h I__4833 (
            .O(N__22090),
            .I(N__22087));
    Span4Mux_s3_v I__4832 (
            .O(N__22087),
            .I(N__22084));
    Odrv4 I__4831 (
            .O(N__22084),
            .I(\sb_translator_1.N_729 ));
    InMux I__4830 (
            .O(N__22081),
            .I(N__22078));
    LocalMux I__4829 (
            .O(N__22078),
            .I(\sb_translator_1.N_712 ));
    InMux I__4828 (
            .O(N__22075),
            .I(N__22067));
    CascadeMux I__4827 (
            .O(N__22074),
            .I(N__22054));
    InMux I__4826 (
            .O(N__22073),
            .I(N__22039));
    InMux I__4825 (
            .O(N__22072),
            .I(N__22036));
    InMux I__4824 (
            .O(N__22071),
            .I(N__22031));
    InMux I__4823 (
            .O(N__22070),
            .I(N__22031));
    LocalMux I__4822 (
            .O(N__22067),
            .I(N__22028));
    InMux I__4821 (
            .O(N__22066),
            .I(N__22025));
    InMux I__4820 (
            .O(N__22065),
            .I(N__22018));
    InMux I__4819 (
            .O(N__22064),
            .I(N__22018));
    InMux I__4818 (
            .O(N__22063),
            .I(N__22018));
    InMux I__4817 (
            .O(N__22062),
            .I(N__22010));
    InMux I__4816 (
            .O(N__22061),
            .I(N__21998));
    InMux I__4815 (
            .O(N__22060),
            .I(N__21998));
    InMux I__4814 (
            .O(N__22059),
            .I(N__21998));
    InMux I__4813 (
            .O(N__22058),
            .I(N__21998));
    InMux I__4812 (
            .O(N__22057),
            .I(N__21998));
    InMux I__4811 (
            .O(N__22054),
            .I(N__21984));
    InMux I__4810 (
            .O(N__22053),
            .I(N__21984));
    InMux I__4809 (
            .O(N__22052),
            .I(N__21977));
    InMux I__4808 (
            .O(N__22051),
            .I(N__21977));
    InMux I__4807 (
            .O(N__22050),
            .I(N__21977));
    InMux I__4806 (
            .O(N__22049),
            .I(N__21966));
    InMux I__4805 (
            .O(N__22048),
            .I(N__21966));
    InMux I__4804 (
            .O(N__22047),
            .I(N__21966));
    InMux I__4803 (
            .O(N__22046),
            .I(N__21966));
    InMux I__4802 (
            .O(N__22045),
            .I(N__21966));
    InMux I__4801 (
            .O(N__22044),
            .I(N__21959));
    InMux I__4800 (
            .O(N__22043),
            .I(N__21959));
    InMux I__4799 (
            .O(N__22042),
            .I(N__21959));
    LocalMux I__4798 (
            .O(N__22039),
            .I(N__21956));
    LocalMux I__4797 (
            .O(N__22036),
            .I(N__21945));
    LocalMux I__4796 (
            .O(N__22031),
            .I(N__21945));
    Span4Mux_v I__4795 (
            .O(N__22028),
            .I(N__21945));
    LocalMux I__4794 (
            .O(N__22025),
            .I(N__21945));
    LocalMux I__4793 (
            .O(N__22018),
            .I(N__21945));
    InMux I__4792 (
            .O(N__22017),
            .I(N__21934));
    InMux I__4791 (
            .O(N__22016),
            .I(N__21934));
    InMux I__4790 (
            .O(N__22015),
            .I(N__21934));
    InMux I__4789 (
            .O(N__22014),
            .I(N__21934));
    InMux I__4788 (
            .O(N__22013),
            .I(N__21934));
    LocalMux I__4787 (
            .O(N__22010),
            .I(N__21931));
    InMux I__4786 (
            .O(N__22009),
            .I(N__21928));
    LocalMux I__4785 (
            .O(N__21998),
            .I(N__21925));
    InMux I__4784 (
            .O(N__21997),
            .I(N__21922));
    InMux I__4783 (
            .O(N__21996),
            .I(N__21905));
    InMux I__4782 (
            .O(N__21995),
            .I(N__21905));
    InMux I__4781 (
            .O(N__21994),
            .I(N__21905));
    InMux I__4780 (
            .O(N__21993),
            .I(N__21905));
    InMux I__4779 (
            .O(N__21992),
            .I(N__21905));
    InMux I__4778 (
            .O(N__21991),
            .I(N__21905));
    InMux I__4777 (
            .O(N__21990),
            .I(N__21905));
    InMux I__4776 (
            .O(N__21989),
            .I(N__21905));
    LocalMux I__4775 (
            .O(N__21984),
            .I(N__21898));
    LocalMux I__4774 (
            .O(N__21977),
            .I(N__21898));
    LocalMux I__4773 (
            .O(N__21966),
            .I(N__21898));
    LocalMux I__4772 (
            .O(N__21959),
            .I(N__21891));
    Span4Mux_v I__4771 (
            .O(N__21956),
            .I(N__21891));
    Span4Mux_v I__4770 (
            .O(N__21945),
            .I(N__21891));
    LocalMux I__4769 (
            .O(N__21934),
            .I(N__21884));
    Span4Mux_v I__4768 (
            .O(N__21931),
            .I(N__21884));
    LocalMux I__4767 (
            .O(N__21928),
            .I(N__21884));
    Span4Mux_v I__4766 (
            .O(N__21925),
            .I(N__21881));
    LocalMux I__4765 (
            .O(N__21922),
            .I(N__21878));
    LocalMux I__4764 (
            .O(N__21905),
            .I(N__21871));
    Span4Mux_v I__4763 (
            .O(N__21898),
            .I(N__21871));
    Span4Mux_h I__4762 (
            .O(N__21891),
            .I(N__21871));
    Span4Mux_v I__4761 (
            .O(N__21884),
            .I(N__21866));
    Span4Mux_h I__4760 (
            .O(N__21881),
            .I(N__21866));
    Span4Mux_v I__4759 (
            .O(N__21878),
            .I(N__21861));
    Span4Mux_h I__4758 (
            .O(N__21871),
            .I(N__21861));
    Odrv4 I__4757 (
            .O(N__21866),
            .I(\sb_translator_1.stateZ0Z_0 ));
    Odrv4 I__4756 (
            .O(N__21861),
            .I(\sb_translator_1.stateZ0Z_0 ));
    InMux I__4755 (
            .O(N__21856),
            .I(N__21852));
    InMux I__4754 (
            .O(N__21855),
            .I(N__21849));
    LocalMux I__4753 (
            .O(N__21852),
            .I(N__21844));
    LocalMux I__4752 (
            .O(N__21849),
            .I(N__21844));
    Span4Mux_v I__4751 (
            .O(N__21844),
            .I(N__21841));
    Span4Mux_h I__4750 (
            .O(N__21841),
            .I(N__21838));
    Odrv4 I__4749 (
            .O(N__21838),
            .I(\sb_translator_1.state_RNIOCIR9Z0Z_5 ));
    InMux I__4748 (
            .O(N__21835),
            .I(N__21832));
    LocalMux I__4747 (
            .O(N__21832),
            .I(\sb_translator_1.state56_a_5_4 ));
    InMux I__4746 (
            .O(N__21829),
            .I(N__21826));
    LocalMux I__4745 (
            .O(N__21826),
            .I(\sb_translator_1.state56_a_5_10 ));
    CascadeMux I__4744 (
            .O(N__21823),
            .I(N__21820));
    InMux I__4743 (
            .O(N__21820),
            .I(N__21817));
    LocalMux I__4742 (
            .O(N__21817),
            .I(\sb_translator_1.state56_a_5_3 ));
    InMux I__4741 (
            .O(N__21814),
            .I(N__21811));
    LocalMux I__4740 (
            .O(N__21811),
            .I(\sb_translator_1.state56_a_5_16 ));
    InMux I__4739 (
            .O(N__21808),
            .I(N__21805));
    LocalMux I__4738 (
            .O(N__21805),
            .I(N__21802));
    Span4Mux_h I__4737 (
            .O(N__21802),
            .I(N__21799));
    Odrv4 I__4736 (
            .O(N__21799),
            .I(demux_data_in_111));
    InMux I__4735 (
            .O(N__21796),
            .I(N__21793));
    LocalMux I__4734 (
            .O(N__21793),
            .I(N__21790));
    Span4Mux_h I__4733 (
            .O(N__21790),
            .I(N__21787));
    Span4Mux_v I__4732 (
            .O(N__21787),
            .I(N__21784));
    Span4Mux_v I__4731 (
            .O(N__21784),
            .I(N__21781));
    Odrv4 I__4730 (
            .O(N__21781),
            .I(demux_data_in_39));
    InMux I__4729 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__4728 (
            .O(N__21775),
            .I(N__21772));
    Span4Mux_h I__4727 (
            .O(N__21772),
            .I(N__21769));
    Span4Mux_v I__4726 (
            .O(N__21769),
            .I(N__21766));
    Odrv4 I__4725 (
            .O(N__21766),
            .I(demux_data_in_95));
    CascadeMux I__4724 (
            .O(N__21763),
            .I(\demux.N_417_i_0_o2Z0Z_0_cascade_ ));
    InMux I__4723 (
            .O(N__21760),
            .I(N__21757));
    LocalMux I__4722 (
            .O(N__21757),
            .I(\demux.N_417_i_0_o2Z0Z_1 ));
    InMux I__4721 (
            .O(N__21754),
            .I(N__21751));
    LocalMux I__4720 (
            .O(N__21751),
            .I(N__21748));
    Span4Mux_v I__4719 (
            .O(N__21748),
            .I(N__21745));
    Span4Mux_h I__4718 (
            .O(N__21745),
            .I(N__21742));
    Odrv4 I__4717 (
            .O(N__21742),
            .I(demux_data_in_47));
    CascadeMux I__4716 (
            .O(N__21739),
            .I(N__21736));
    InMux I__4715 (
            .O(N__21736),
            .I(N__21733));
    LocalMux I__4714 (
            .O(N__21733),
            .I(\demux.N_417_i_0_a3Z0Z_4 ));
    InMux I__4713 (
            .O(N__21730),
            .I(N__21727));
    LocalMux I__4712 (
            .O(N__21727),
            .I(N__21724));
    Span4Mux_h I__4711 (
            .O(N__21724),
            .I(N__21721));
    Odrv4 I__4710 (
            .O(N__21721),
            .I(demux_data_in_109));
    InMux I__4709 (
            .O(N__21718),
            .I(N__21715));
    LocalMux I__4708 (
            .O(N__21715),
            .I(N__21712));
    Span4Mux_h I__4707 (
            .O(N__21712),
            .I(N__21709));
    Span4Mux_v I__4706 (
            .O(N__21709),
            .I(N__21706));
    Span4Mux_v I__4705 (
            .O(N__21706),
            .I(N__21703));
    Odrv4 I__4704 (
            .O(N__21703),
            .I(demux_data_in_37));
    InMux I__4703 (
            .O(N__21700),
            .I(N__21697));
    LocalMux I__4702 (
            .O(N__21697),
            .I(N__21694));
    Span4Mux_h I__4701 (
            .O(N__21694),
            .I(N__21691));
    Span4Mux_v I__4700 (
            .O(N__21691),
            .I(N__21688));
    Odrv4 I__4699 (
            .O(N__21688),
            .I(demux_data_in_93));
    CascadeMux I__4698 (
            .O(N__21685),
            .I(\demux.N_419_i_0_o2Z0Z_0_cascade_ ));
    InMux I__4697 (
            .O(N__21682),
            .I(N__21679));
    LocalMux I__4696 (
            .O(N__21679),
            .I(N__21676));
    Span4Mux_v I__4695 (
            .O(N__21676),
            .I(N__21673));
    Span4Mux_h I__4694 (
            .O(N__21673),
            .I(N__21670));
    Odrv4 I__4693 (
            .O(N__21670),
            .I(demux_data_in_45));
    CascadeMux I__4692 (
            .O(N__21667),
            .I(\demux.N_419_i_0_o2Z0Z_2_cascade_ ));
    InMux I__4691 (
            .O(N__21664),
            .I(N__21661));
    LocalMux I__4690 (
            .O(N__21661),
            .I(N__21658));
    Odrv4 I__4689 (
            .O(N__21658),
            .I(demux_data_in_13));
    InMux I__4688 (
            .O(N__21655),
            .I(N__21652));
    LocalMux I__4687 (
            .O(N__21652),
            .I(\demux.N_419_i_0_a3Z0Z_5 ));
    CascadeMux I__4686 (
            .O(N__21649),
            .I(N__21646));
    InMux I__4685 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__4684 (
            .O(N__21643),
            .I(N__21640));
    Span4Mux_s3_v I__4683 (
            .O(N__21640),
            .I(N__21637));
    Span4Mux_h I__4682 (
            .O(N__21637),
            .I(N__21634));
    Odrv4 I__4681 (
            .O(N__21634),
            .I(demux_data_in_69));
    InMux I__4680 (
            .O(N__21631),
            .I(N__21628));
    LocalMux I__4679 (
            .O(N__21628),
            .I(\demux.N_419_i_0_a3Z0Z_7 ));
    InMux I__4678 (
            .O(N__21625),
            .I(N__21622));
    LocalMux I__4677 (
            .O(N__21622),
            .I(\demux.N_419_i_0_o2Z0Z_8 ));
    InMux I__4676 (
            .O(N__21619),
            .I(N__21616));
    LocalMux I__4675 (
            .O(N__21616),
            .I(N__21611));
    InMux I__4674 (
            .O(N__21615),
            .I(N__21608));
    InMux I__4673 (
            .O(N__21614),
            .I(N__21605));
    Span4Mux_h I__4672 (
            .O(N__21611),
            .I(N__21601));
    LocalMux I__4671 (
            .O(N__21608),
            .I(N__21598));
    LocalMux I__4670 (
            .O(N__21605),
            .I(N__21595));
    InMux I__4669 (
            .O(N__21604),
            .I(N__21592));
    Odrv4 I__4668 (
            .O(N__21601),
            .I(\demux.N_422_i_0_o2Z0Z_9 ));
    Odrv4 I__4667 (
            .O(N__21598),
            .I(\demux.N_422_i_0_o2Z0Z_9 ));
    Odrv4 I__4666 (
            .O(N__21595),
            .I(\demux.N_422_i_0_o2Z0Z_9 ));
    LocalMux I__4665 (
            .O(N__21592),
            .I(\demux.N_422_i_0_o2Z0Z_9 ));
    CascadeMux I__4664 (
            .O(N__21583),
            .I(N__21580));
    InMux I__4663 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__4662 (
            .O(N__21577),
            .I(N__21571));
    CascadeMux I__4661 (
            .O(N__21576),
            .I(N__21568));
    CascadeMux I__4660 (
            .O(N__21575),
            .I(N__21565));
    CascadeMux I__4659 (
            .O(N__21574),
            .I(N__21562));
    Span4Mux_h I__4658 (
            .O(N__21571),
            .I(N__21559));
    InMux I__4657 (
            .O(N__21568),
            .I(N__21556));
    InMux I__4656 (
            .O(N__21565),
            .I(N__21553));
    InMux I__4655 (
            .O(N__21562),
            .I(N__21550));
    Odrv4 I__4654 (
            .O(N__21559),
            .I(\demux.N_422_i_0_aZ0Z3 ));
    LocalMux I__4653 (
            .O(N__21556),
            .I(\demux.N_422_i_0_aZ0Z3 ));
    LocalMux I__4652 (
            .O(N__21553),
            .I(\demux.N_422_i_0_aZ0Z3 ));
    LocalMux I__4651 (
            .O(N__21550),
            .I(\demux.N_422_i_0_aZ0Z3 ));
    InMux I__4650 (
            .O(N__21541),
            .I(N__21535));
    InMux I__4649 (
            .O(N__21540),
            .I(N__21532));
    InMux I__4648 (
            .O(N__21539),
            .I(N__21529));
    InMux I__4647 (
            .O(N__21538),
            .I(N__21526));
    LocalMux I__4646 (
            .O(N__21535),
            .I(\demux.N_422_i_0_o2Z0Z_7 ));
    LocalMux I__4645 (
            .O(N__21532),
            .I(\demux.N_422_i_0_o2Z0Z_7 ));
    LocalMux I__4644 (
            .O(N__21529),
            .I(\demux.N_422_i_0_o2Z0Z_7 ));
    LocalMux I__4643 (
            .O(N__21526),
            .I(\demux.N_422_i_0_o2Z0Z_7 ));
    CEMux I__4642 (
            .O(N__21517),
            .I(N__21513));
    CEMux I__4641 (
            .O(N__21516),
            .I(N__21510));
    LocalMux I__4640 (
            .O(N__21513),
            .I(N__21507));
    LocalMux I__4639 (
            .O(N__21510),
            .I(N__21504));
    Span4Mux_v I__4638 (
            .O(N__21507),
            .I(N__21500));
    Span4Mux_v I__4637 (
            .O(N__21504),
            .I(N__21497));
    CEMux I__4636 (
            .O(N__21503),
            .I(N__21494));
    Span4Mux_h I__4635 (
            .O(N__21500),
            .I(N__21491));
    Span4Mux_v I__4634 (
            .O(N__21497),
            .I(N__21488));
    LocalMux I__4633 (
            .O(N__21494),
            .I(N__21485));
    Span4Mux_v I__4632 (
            .O(N__21491),
            .I(N__21482));
    Sp12to4 I__4631 (
            .O(N__21488),
            .I(N__21479));
    Span12Mux_s11_v I__4630 (
            .O(N__21485),
            .I(N__21476));
    Odrv4 I__4629 (
            .O(N__21482),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1 ));
    Odrv12 I__4628 (
            .O(N__21479),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1 ));
    Odrv12 I__4627 (
            .O(N__21476),
            .I(\sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1 ));
    InMux I__4626 (
            .O(N__21469),
            .I(N__21466));
    LocalMux I__4625 (
            .O(N__21466),
            .I(N__21463));
    Span4Mux_v I__4624 (
            .O(N__21463),
            .I(N__21460));
    Odrv4 I__4623 (
            .O(N__21460),
            .I(mosi_data_out_16));
    InMux I__4622 (
            .O(N__21457),
            .I(N__21454));
    LocalMux I__4621 (
            .O(N__21454),
            .I(N__21451));
    Span4Mux_h I__4620 (
            .O(N__21451),
            .I(N__21448));
    Span4Mux_v I__4619 (
            .O(N__21448),
            .I(N__21443));
    InMux I__4618 (
            .O(N__21447),
            .I(N__21440));
    InMux I__4617 (
            .O(N__21446),
            .I(N__21437));
    Odrv4 I__4616 (
            .O(N__21443),
            .I(\sb_translator_1.cntZ0Z_8 ));
    LocalMux I__4615 (
            .O(N__21440),
            .I(\sb_translator_1.cntZ0Z_8 ));
    LocalMux I__4614 (
            .O(N__21437),
            .I(\sb_translator_1.cntZ0Z_8 ));
    InMux I__4613 (
            .O(N__21430),
            .I(N__21427));
    LocalMux I__4612 (
            .O(N__21427),
            .I(N__21424));
    Span4Mux_h I__4611 (
            .O(N__21424),
            .I(N__21421));
    Odrv4 I__4610 (
            .O(N__21421),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_8 ));
    CascadeMux I__4609 (
            .O(N__21418),
            .I(N__21413));
    CascadeMux I__4608 (
            .O(N__21417),
            .I(N__21410));
    InMux I__4607 (
            .O(N__21416),
            .I(N__21406));
    InMux I__4606 (
            .O(N__21413),
            .I(N__21399));
    InMux I__4605 (
            .O(N__21410),
            .I(N__21399));
    InMux I__4604 (
            .O(N__21409),
            .I(N__21399));
    LocalMux I__4603 (
            .O(N__21406),
            .I(N__21395));
    LocalMux I__4602 (
            .O(N__21399),
            .I(N__21392));
    CascadeMux I__4601 (
            .O(N__21398),
            .I(N__21388));
    Span4Mux_v I__4600 (
            .O(N__21395),
            .I(N__21384));
    Span4Mux_h I__4599 (
            .O(N__21392),
            .I(N__21381));
    InMux I__4598 (
            .O(N__21391),
            .I(N__21378));
    InMux I__4597 (
            .O(N__21388),
            .I(N__21373));
    InMux I__4596 (
            .O(N__21387),
            .I(N__21373));
    Odrv4 I__4595 (
            .O(N__21384),
            .I(\sb_translator_1.cnt_ledsZ0Z_12 ));
    Odrv4 I__4594 (
            .O(N__21381),
            .I(\sb_translator_1.cnt_ledsZ0Z_12 ));
    LocalMux I__4593 (
            .O(N__21378),
            .I(\sb_translator_1.cnt_ledsZ0Z_12 ));
    LocalMux I__4592 (
            .O(N__21373),
            .I(\sb_translator_1.cnt_ledsZ0Z_12 ));
    CascadeMux I__4591 (
            .O(N__21364),
            .I(N__21357));
    InMux I__4590 (
            .O(N__21363),
            .I(N__21353));
    InMux I__4589 (
            .O(N__21362),
            .I(N__21345));
    InMux I__4588 (
            .O(N__21361),
            .I(N__21345));
    InMux I__4587 (
            .O(N__21360),
            .I(N__21345));
    InMux I__4586 (
            .O(N__21357),
            .I(N__21340));
    InMux I__4585 (
            .O(N__21356),
            .I(N__21340));
    LocalMux I__4584 (
            .O(N__21353),
            .I(N__21337));
    InMux I__4583 (
            .O(N__21352),
            .I(N__21334));
    LocalMux I__4582 (
            .O(N__21345),
            .I(N__21331));
    LocalMux I__4581 (
            .O(N__21340),
            .I(N__21328));
    Span4Mux_v I__4580 (
            .O(N__21337),
            .I(N__21325));
    LocalMux I__4579 (
            .O(N__21334),
            .I(N__21318));
    Span4Mux_v I__4578 (
            .O(N__21331),
            .I(N__21318));
    Span4Mux_v I__4577 (
            .O(N__21328),
            .I(N__21318));
    Odrv4 I__4576 (
            .O(N__21325),
            .I(\sb_translator_1.cnt_ledsZ0Z_9 ));
    Odrv4 I__4575 (
            .O(N__21318),
            .I(\sb_translator_1.cnt_ledsZ0Z_9 ));
    InMux I__4574 (
            .O(N__21313),
            .I(N__21307));
    InMux I__4573 (
            .O(N__21312),
            .I(N__21300));
    InMux I__4572 (
            .O(N__21311),
            .I(N__21300));
    InMux I__4571 (
            .O(N__21310),
            .I(N__21300));
    LocalMux I__4570 (
            .O(N__21307),
            .I(N__21297));
    LocalMux I__4569 (
            .O(N__21300),
            .I(N__21294));
    Span4Mux_h I__4568 (
            .O(N__21297),
            .I(N__21289));
    Span4Mux_v I__4567 (
            .O(N__21294),
            .I(N__21289));
    Span4Mux_h I__4566 (
            .O(N__21289),
            .I(N__21286));
    Odrv4 I__4565 (
            .O(N__21286),
            .I(\sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9 ));
    CascadeMux I__4564 (
            .O(N__21283),
            .I(N__21280));
    InMux I__4563 (
            .O(N__21280),
            .I(N__21277));
    LocalMux I__4562 (
            .O(N__21277),
            .I(N__21274));
    Span12Mux_v I__4561 (
            .O(N__21274),
            .I(N__21271));
    Odrv12 I__4560 (
            .O(N__21271),
            .I(demux_data_in_26));
    InMux I__4559 (
            .O(N__21268),
            .I(N__21265));
    LocalMux I__4558 (
            .O(N__21265),
            .I(N__21262));
    Odrv4 I__4557 (
            .O(N__21262),
            .I(\demux.N_422_i_0_a3Z0Z_7 ));
    InMux I__4556 (
            .O(N__21259),
            .I(N__21256));
    LocalMux I__4555 (
            .O(N__21256),
            .I(N__21253));
    Span4Mux_v I__4554 (
            .O(N__21253),
            .I(N__21250));
    Odrv4 I__4553 (
            .O(N__21250),
            .I(demux_data_in_15));
    InMux I__4552 (
            .O(N__21247),
            .I(N__21244));
    LocalMux I__4551 (
            .O(N__21244),
            .I(N__21241));
    Span4Mux_h I__4550 (
            .O(N__21241),
            .I(N__21238));
    Span4Mux_v I__4549 (
            .O(N__21238),
            .I(N__21235));
    Span4Mux_v I__4548 (
            .O(N__21235),
            .I(N__21232));
    Odrv4 I__4547 (
            .O(N__21232),
            .I(demux_data_in_25));
    InMux I__4546 (
            .O(N__21229),
            .I(N__21226));
    LocalMux I__4545 (
            .O(N__21226),
            .I(N__21223));
    Span4Mux_h I__4544 (
            .O(N__21223),
            .I(N__21220));
    Odrv4 I__4543 (
            .O(N__21220),
            .I(demux_data_in_17));
    CascadeMux I__4542 (
            .O(N__21217),
            .I(N__21214));
    InMux I__4541 (
            .O(N__21214),
            .I(N__21211));
    LocalMux I__4540 (
            .O(N__21211),
            .I(N__21208));
    Span4Mux_h I__4539 (
            .O(N__21208),
            .I(N__21205));
    Odrv4 I__4538 (
            .O(N__21205),
            .I(demux_data_in_97));
    InMux I__4537 (
            .O(N__21202),
            .I(N__21199));
    LocalMux I__4536 (
            .O(N__21199),
            .I(N__21196));
    Span4Mux_h I__4535 (
            .O(N__21196),
            .I(N__21193));
    Span4Mux_h I__4534 (
            .O(N__21193),
            .I(N__21190));
    Odrv4 I__4533 (
            .O(N__21190),
            .I(demux_data_in_65));
    CascadeMux I__4532 (
            .O(N__21187),
            .I(\demux.N_423_i_0_o2Z0Z_4_cascade_ ));
    InMux I__4531 (
            .O(N__21184),
            .I(N__21181));
    LocalMux I__4530 (
            .O(N__21181),
            .I(\demux.N_423_i_0_a3Z0Z_7 ));
    InMux I__4529 (
            .O(N__21178),
            .I(N__21175));
    LocalMux I__4528 (
            .O(N__21175),
            .I(N__21172));
    Span4Mux_h I__4527 (
            .O(N__21172),
            .I(N__21169));
    Span4Mux_v I__4526 (
            .O(N__21169),
            .I(N__21166));
    Odrv4 I__4525 (
            .O(N__21166),
            .I(demux_data_in_41));
    CascadeMux I__4524 (
            .O(N__21163),
            .I(\demux.N_423_i_0_o2Z0Z_8_cascade_ ));
    InMux I__4523 (
            .O(N__21160),
            .I(N__21157));
    LocalMux I__4522 (
            .O(N__21157),
            .I(\demux.N_423_i_0_o2Z0Z_2 ));
    InMux I__4521 (
            .O(N__21154),
            .I(N__21151));
    LocalMux I__4520 (
            .O(N__21151),
            .I(\demux.N_418_i_0_o2Z0Z_4 ));
    InMux I__4519 (
            .O(N__21148),
            .I(N__21145));
    LocalMux I__4518 (
            .O(N__21145),
            .I(N__21142));
    Span4Mux_v I__4517 (
            .O(N__21142),
            .I(N__21139));
    Span4Mux_h I__4516 (
            .O(N__21139),
            .I(N__21136));
    Odrv4 I__4515 (
            .O(N__21136),
            .I(demux_data_in_78));
    CascadeMux I__4514 (
            .O(N__21133),
            .I(\demux.N_884_cascade_ ));
    InMux I__4513 (
            .O(N__21130),
            .I(N__21127));
    LocalMux I__4512 (
            .O(N__21127),
            .I(N__21124));
    Span4Mux_v I__4511 (
            .O(N__21124),
            .I(N__21121));
    Span4Mux_h I__4510 (
            .O(N__21121),
            .I(N__21118));
    Odrv4 I__4509 (
            .O(N__21118),
            .I(demux_data_in_27));
    InMux I__4508 (
            .O(N__21115),
            .I(N__21112));
    LocalMux I__4507 (
            .O(N__21112),
            .I(N__21109));
    Span4Mux_h I__4506 (
            .O(N__21109),
            .I(N__21106));
    Span4Mux_v I__4505 (
            .O(N__21106),
            .I(N__21103));
    Odrv4 I__4504 (
            .O(N__21103),
            .I(demux_data_in_19));
    CascadeMux I__4503 (
            .O(N__21100),
            .I(N__21097));
    InMux I__4502 (
            .O(N__21097),
            .I(N__21094));
    LocalMux I__4501 (
            .O(N__21094),
            .I(N__21091));
    Odrv4 I__4500 (
            .O(N__21091),
            .I(demux_data_in_99));
    InMux I__4499 (
            .O(N__21088),
            .I(N__21085));
    LocalMux I__4498 (
            .O(N__21085),
            .I(N__21082));
    Span4Mux_v I__4497 (
            .O(N__21082),
            .I(N__21079));
    Span4Mux_h I__4496 (
            .O(N__21079),
            .I(N__21076));
    Odrv4 I__4495 (
            .O(N__21076),
            .I(demux_data_in_75));
    InMux I__4494 (
            .O(N__21073),
            .I(N__21064));
    InMux I__4493 (
            .O(N__21072),
            .I(N__21064));
    CascadeMux I__4492 (
            .O(N__21071),
            .I(N__21061));
    CascadeMux I__4491 (
            .O(N__21070),
            .I(N__21056));
    CascadeMux I__4490 (
            .O(N__21069),
            .I(N__21053));
    LocalMux I__4489 (
            .O(N__21064),
            .I(N__21049));
    InMux I__4488 (
            .O(N__21061),
            .I(N__21042));
    InMux I__4487 (
            .O(N__21060),
            .I(N__21042));
    InMux I__4486 (
            .O(N__21059),
            .I(N__21042));
    InMux I__4485 (
            .O(N__21056),
            .I(N__21035));
    InMux I__4484 (
            .O(N__21053),
            .I(N__21035));
    InMux I__4483 (
            .O(N__21052),
            .I(N__21035));
    Span4Mux_h I__4482 (
            .O(N__21049),
            .I(N__21030));
    LocalMux I__4481 (
            .O(N__21042),
            .I(N__21030));
    LocalMux I__4480 (
            .O(N__21035),
            .I(\demux.N_424_i_0_a2Z0Z_0 ));
    Odrv4 I__4479 (
            .O(N__21030),
            .I(\demux.N_424_i_0_a2Z0Z_0 ));
    CascadeMux I__4478 (
            .O(N__21025),
            .I(\demux.N_421_i_0_o2Z0Z_4_cascade_ ));
    InMux I__4477 (
            .O(N__21022),
            .I(N__21019));
    LocalMux I__4476 (
            .O(N__21019),
            .I(\demux.N_421_i_0_a3Z0Z_7 ));
    InMux I__4475 (
            .O(N__21016),
            .I(N__21013));
    LocalMux I__4474 (
            .O(N__21013),
            .I(N__21010));
    Span4Mux_h I__4473 (
            .O(N__21010),
            .I(N__21007));
    Odrv4 I__4472 (
            .O(N__21007),
            .I(demux_data_in_11));
    CascadeMux I__4471 (
            .O(N__21004),
            .I(\demux.N_421_i_0_o2Z0Z_8_cascade_ ));
    InMux I__4470 (
            .O(N__21001),
            .I(N__20998));
    LocalMux I__4469 (
            .O(N__20998),
            .I(\demux.N_421_i_0_o2Z0Z_2 ));
    InMux I__4468 (
            .O(N__20995),
            .I(N__20991));
    InMux I__4467 (
            .O(N__20994),
            .I(N__20987));
    LocalMux I__4466 (
            .O(N__20991),
            .I(N__20984));
    InMux I__4465 (
            .O(N__20990),
            .I(N__20981));
    LocalMux I__4464 (
            .O(N__20987),
            .I(N__20977));
    Span4Mux_h I__4463 (
            .O(N__20984),
            .I(N__20972));
    LocalMux I__4462 (
            .O(N__20981),
            .I(N__20972));
    InMux I__4461 (
            .O(N__20980),
            .I(N__20969));
    Odrv4 I__4460 (
            .O(N__20977),
            .I(\demux.N_422_i_0_o2Z0Z_8 ));
    Odrv4 I__4459 (
            .O(N__20972),
            .I(\demux.N_422_i_0_o2Z0Z_8 ));
    LocalMux I__4458 (
            .O(N__20969),
            .I(\demux.N_422_i_0_o2Z0Z_8 ));
    CascadeMux I__4457 (
            .O(N__20962),
            .I(N__20958));
    InMux I__4456 (
            .O(N__20961),
            .I(N__20953));
    InMux I__4455 (
            .O(N__20958),
            .I(N__20953));
    LocalMux I__4454 (
            .O(N__20953),
            .I(N__20950));
    Span4Mux_v I__4453 (
            .O(N__20950),
            .I(N__20943));
    InMux I__4452 (
            .O(N__20949),
            .I(N__20940));
    InMux I__4451 (
            .O(N__20948),
            .I(N__20937));
    InMux I__4450 (
            .O(N__20947),
            .I(N__20932));
    InMux I__4449 (
            .O(N__20946),
            .I(N__20932));
    Span4Mux_h I__4448 (
            .O(N__20943),
            .I(N__20929));
    LocalMux I__4447 (
            .O(N__20940),
            .I(\sb_translator_1.num_ledsZ0Z_15 ));
    LocalMux I__4446 (
            .O(N__20937),
            .I(\sb_translator_1.num_ledsZ0Z_15 ));
    LocalMux I__4445 (
            .O(N__20932),
            .I(\sb_translator_1.num_ledsZ0Z_15 ));
    Odrv4 I__4444 (
            .O(N__20929),
            .I(\sb_translator_1.num_ledsZ0Z_15 ));
    CascadeMux I__4443 (
            .O(N__20920),
            .I(N__20917));
    InMux I__4442 (
            .O(N__20917),
            .I(N__20913));
    InMux I__4441 (
            .O(N__20916),
            .I(N__20910));
    LocalMux I__4440 (
            .O(N__20913),
            .I(\sb_translator_1.cnt_leds_i_16 ));
    LocalMux I__4439 (
            .O(N__20910),
            .I(\sb_translator_1.cnt_leds_i_16 ));
    InMux I__4438 (
            .O(N__20905),
            .I(N__20900));
    InMux I__4437 (
            .O(N__20904),
            .I(N__20895));
    InMux I__4436 (
            .O(N__20903),
            .I(N__20895));
    LocalMux I__4435 (
            .O(N__20900),
            .I(\sb_translator_1.cnt_ledsZ0Z_15 ));
    LocalMux I__4434 (
            .O(N__20895),
            .I(\sb_translator_1.cnt_ledsZ0Z_15 ));
    CascadeMux I__4433 (
            .O(N__20890),
            .I(N__20887));
    InMux I__4432 (
            .O(N__20887),
            .I(N__20884));
    LocalMux I__4431 (
            .O(N__20884),
            .I(N__20881));
    Odrv4 I__4430 (
            .O(N__20881),
            .I(\sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15 ));
    InMux I__4429 (
            .O(N__20878),
            .I(N__20871));
    InMux I__4428 (
            .O(N__20877),
            .I(N__20871));
    CascadeMux I__4427 (
            .O(N__20876),
            .I(N__20867));
    LocalMux I__4426 (
            .O(N__20871),
            .I(N__20862));
    InMux I__4425 (
            .O(N__20870),
            .I(N__20857));
    InMux I__4424 (
            .O(N__20867),
            .I(N__20857));
    InMux I__4423 (
            .O(N__20866),
            .I(N__20852));
    InMux I__4422 (
            .O(N__20865),
            .I(N__20852));
    Span4Mux_v I__4421 (
            .O(N__20862),
            .I(N__20849));
    LocalMux I__4420 (
            .O(N__20857),
            .I(\sb_translator_1.num_ledsZ0Z_12 ));
    LocalMux I__4419 (
            .O(N__20852),
            .I(\sb_translator_1.num_ledsZ0Z_12 ));
    Odrv4 I__4418 (
            .O(N__20849),
            .I(\sb_translator_1.num_ledsZ0Z_12 ));
    InMux I__4417 (
            .O(N__20842),
            .I(N__20837));
    InMux I__4416 (
            .O(N__20841),
            .I(N__20832));
    InMux I__4415 (
            .O(N__20840),
            .I(N__20832));
    LocalMux I__4414 (
            .O(N__20837),
            .I(\sb_translator_1.cnt_ledsZ0Z_13 ));
    LocalMux I__4413 (
            .O(N__20832),
            .I(\sb_translator_1.cnt_ledsZ0Z_13 ));
    InMux I__4412 (
            .O(N__20827),
            .I(N__20824));
    LocalMux I__4411 (
            .O(N__20824),
            .I(N__20821));
    Span4Mux_s3_v I__4410 (
            .O(N__20821),
            .I(N__20818));
    Odrv4 I__4409 (
            .O(N__20818),
            .I(\sb_translator_1.cnt_leds_RNI15HTZ0Z_13 ));
    InMux I__4408 (
            .O(N__20815),
            .I(N__20803));
    InMux I__4407 (
            .O(N__20814),
            .I(N__20803));
    InMux I__4406 (
            .O(N__20813),
            .I(N__20803));
    InMux I__4405 (
            .O(N__20812),
            .I(N__20803));
    LocalMux I__4404 (
            .O(N__20803),
            .I(N__20799));
    CascadeMux I__4403 (
            .O(N__20802),
            .I(N__20795));
    Span4Mux_h I__4402 (
            .O(N__20799),
            .I(N__20792));
    InMux I__4401 (
            .O(N__20798),
            .I(N__20787));
    InMux I__4400 (
            .O(N__20795),
            .I(N__20787));
    Odrv4 I__4399 (
            .O(N__20792),
            .I(\sb_translator_1.num_ledsZ0Z_14 ));
    LocalMux I__4398 (
            .O(N__20787),
            .I(\sb_translator_1.num_ledsZ0Z_14 ));
    CascadeMux I__4397 (
            .O(N__20782),
            .I(N__20777));
    InMux I__4396 (
            .O(N__20781),
            .I(N__20766));
    InMux I__4395 (
            .O(N__20780),
            .I(N__20766));
    InMux I__4394 (
            .O(N__20777),
            .I(N__20766));
    InMux I__4393 (
            .O(N__20776),
            .I(N__20766));
    CascadeMux I__4392 (
            .O(N__20775),
            .I(N__20762));
    LocalMux I__4391 (
            .O(N__20766),
            .I(N__20759));
    InMux I__4390 (
            .O(N__20765),
            .I(N__20754));
    InMux I__4389 (
            .O(N__20762),
            .I(N__20754));
    Span4Mux_h I__4388 (
            .O(N__20759),
            .I(N__20751));
    LocalMux I__4387 (
            .O(N__20754),
            .I(\sb_translator_1.num_ledsZ0Z_13 ));
    Odrv4 I__4386 (
            .O(N__20751),
            .I(\sb_translator_1.num_ledsZ0Z_13 ));
    CascadeMux I__4385 (
            .O(N__20746),
            .I(\sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_ ));
    InMux I__4384 (
            .O(N__20743),
            .I(N__20738));
    InMux I__4383 (
            .O(N__20742),
            .I(N__20733));
    InMux I__4382 (
            .O(N__20741),
            .I(N__20733));
    LocalMux I__4381 (
            .O(N__20738),
            .I(\sb_translator_1.cnt_ledsZ0Z_14 ));
    LocalMux I__4380 (
            .O(N__20733),
            .I(\sb_translator_1.cnt_ledsZ0Z_14 ));
    CascadeMux I__4379 (
            .O(N__20728),
            .I(N__20725));
    InMux I__4378 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__4377 (
            .O(N__20722),
            .I(N__20719));
    Odrv4 I__4376 (
            .O(N__20719),
            .I(\sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14 ));
    CascadeMux I__4375 (
            .O(N__20716),
            .I(N__20713));
    InMux I__4374 (
            .O(N__20713),
            .I(N__20710));
    LocalMux I__4373 (
            .O(N__20710),
            .I(N__20707));
    Span12Mux_s11_v I__4372 (
            .O(N__20707),
            .I(N__20704));
    Odrv12 I__4371 (
            .O(N__20704),
            .I(demux_data_in_66));
    InMux I__4370 (
            .O(N__20701),
            .I(N__20698));
    LocalMux I__4369 (
            .O(N__20698),
            .I(N__20695));
    Span4Mux_v I__4368 (
            .O(N__20695),
            .I(N__20692));
    Span4Mux_h I__4367 (
            .O(N__20692),
            .I(N__20689));
    Odrv4 I__4366 (
            .O(N__20689),
            .I(demux_data_in_30));
    CascadeMux I__4365 (
            .O(N__20686),
            .I(N__20683));
    InMux I__4364 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__4363 (
            .O(N__20680),
            .I(N__20677));
    Odrv4 I__4362 (
            .O(N__20677),
            .I(demux_data_in_102));
    InMux I__4361 (
            .O(N__20674),
            .I(N__20671));
    LocalMux I__4360 (
            .O(N__20671),
            .I(N__20668));
    Span4Mux_h I__4359 (
            .O(N__20668),
            .I(N__20665));
    Span4Mux_h I__4358 (
            .O(N__20665),
            .I(N__20662));
    Odrv4 I__4357 (
            .O(N__20662),
            .I(demux_data_in_32));
    CascadeMux I__4356 (
            .O(N__20659),
            .I(N__20656));
    InMux I__4355 (
            .O(N__20656),
            .I(N__20653));
    LocalMux I__4354 (
            .O(N__20653),
            .I(N__20650));
    Span4Mux_h I__4353 (
            .O(N__20650),
            .I(N__20647));
    Odrv4 I__4352 (
            .O(N__20647),
            .I(demux_data_in_104));
    InMux I__4351 (
            .O(N__20644),
            .I(N__20641));
    LocalMux I__4350 (
            .O(N__20641),
            .I(\demux.N_424_i_0_o2_0Z0Z_0 ));
    InMux I__4349 (
            .O(N__20638),
            .I(N__20635));
    LocalMux I__4348 (
            .O(N__20635),
            .I(N__20632));
    Span4Mux_h I__4347 (
            .O(N__20632),
            .I(N__20629));
    Span4Mux_h I__4346 (
            .O(N__20629),
            .I(N__20626));
    Odrv4 I__4345 (
            .O(N__20626),
            .I(demux_data_in_44));
    InMux I__4344 (
            .O(N__20623),
            .I(N__20620));
    LocalMux I__4343 (
            .O(N__20620),
            .I(N__20617));
    Span4Mux_h I__4342 (
            .O(N__20617),
            .I(N__20614));
    Span4Mux_v I__4341 (
            .O(N__20614),
            .I(N__20611));
    Odrv4 I__4340 (
            .O(N__20611),
            .I(demux_data_in_22));
    InMux I__4339 (
            .O(N__20608),
            .I(\sb_translator_1.state56_a_5_cry_12 ));
    InMux I__4338 (
            .O(N__20605),
            .I(\sb_translator_1.state56_a_5_cry_13 ));
    InMux I__4337 (
            .O(N__20602),
            .I(bfn_8_5_0_));
    InMux I__4336 (
            .O(N__20599),
            .I(N__20595));
    InMux I__4335 (
            .O(N__20598),
            .I(N__20592));
    LocalMux I__4334 (
            .O(N__20595),
            .I(\sb_translator_1.cnt_ledsZ0Z_16 ));
    LocalMux I__4333 (
            .O(N__20592),
            .I(\sb_translator_1.cnt_ledsZ0Z_16 ));
    CascadeMux I__4332 (
            .O(N__20587),
            .I(\sb_translator_1.cnt_leds_i_16_cascade_ ));
    InMux I__4331 (
            .O(N__20584),
            .I(N__20581));
    LocalMux I__4330 (
            .O(N__20581),
            .I(N__20578));
    Odrv4 I__4329 (
            .O(N__20578),
            .I(\sb_translator_1.num_leds_RNIOJBMZ0Z_15 ));
    InMux I__4328 (
            .O(N__20575),
            .I(N__20571));
    CascadeMux I__4327 (
            .O(N__20574),
            .I(N__20568));
    LocalMux I__4326 (
            .O(N__20571),
            .I(N__20565));
    InMux I__4325 (
            .O(N__20568),
            .I(N__20562));
    Span4Mux_v I__4324 (
            .O(N__20565),
            .I(N__20557));
    LocalMux I__4323 (
            .O(N__20562),
            .I(N__20557));
    Odrv4 I__4322 (
            .O(N__20557),
            .I(\sb_translator_1.num_leds_RNIU1HTZ0Z_11 ));
    InMux I__4321 (
            .O(N__20554),
            .I(N__20551));
    LocalMux I__4320 (
            .O(N__20551),
            .I(N__20548));
    Odrv4 I__4319 (
            .O(N__20548),
            .I(\sb_translator_1.cnt_leds_RNIV62R1Z0Z_13 ));
    CascadeMux I__4318 (
            .O(N__20545),
            .I(N__20542));
    InMux I__4317 (
            .O(N__20542),
            .I(N__20539));
    LocalMux I__4316 (
            .O(N__20539),
            .I(N__20536));
    Odrv4 I__4315 (
            .O(N__20536),
            .I(\sb_translator_1.cnt_leds_RNI48HTZ0Z_14 ));
    CascadeMux I__4314 (
            .O(N__20533),
            .I(\sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_ ));
    InMux I__4313 (
            .O(N__20530),
            .I(N__20527));
    LocalMux I__4312 (
            .O(N__20527),
            .I(N__20524));
    Odrv4 I__4311 (
            .O(N__20524),
            .I(\sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15 ));
    InMux I__4310 (
            .O(N__20521),
            .I(N__20518));
    LocalMux I__4309 (
            .O(N__20518),
            .I(\sb_translator_1.cnt_leds_RNIHCUTZ0Z_7 ));
    CascadeMux I__4308 (
            .O(N__20515),
            .I(N__20512));
    InMux I__4307 (
            .O(N__20512),
            .I(N__20509));
    LocalMux I__4306 (
            .O(N__20509),
            .I(\sb_translator_1.cnt_leds_RNIN4VEZ0Z_6 ));
    InMux I__4305 (
            .O(N__20506),
            .I(\sb_translator_1.state56_a_5_cry_4 ));
    InMux I__4304 (
            .O(N__20503),
            .I(N__20500));
    LocalMux I__4303 (
            .O(N__20500),
            .I(\sb_translator_1.cnt_leds_RNINIUTZ0Z_8 ));
    CascadeMux I__4302 (
            .O(N__20497),
            .I(N__20494));
    InMux I__4301 (
            .O(N__20494),
            .I(N__20491));
    LocalMux I__4300 (
            .O(N__20491),
            .I(\sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7 ));
    InMux I__4299 (
            .O(N__20488),
            .I(\sb_translator_1.state56_a_5_cry_5 ));
    InMux I__4298 (
            .O(N__20485),
            .I(N__20482));
    LocalMux I__4297 (
            .O(N__20482),
            .I(N__20479));
    Odrv4 I__4296 (
            .O(N__20479),
            .I(\sb_translator_1.num_leds_RNITOUTZ0Z_8 ));
    InMux I__4295 (
            .O(N__20476),
            .I(N__20472));
    CascadeMux I__4294 (
            .O(N__20475),
            .I(N__20469));
    LocalMux I__4293 (
            .O(N__20472),
            .I(N__20466));
    InMux I__4292 (
            .O(N__20469),
            .I(N__20463));
    Span4Mux_v I__4291 (
            .O(N__20466),
            .I(N__20460));
    LocalMux I__4290 (
            .O(N__20463),
            .I(N__20457));
    Odrv4 I__4289 (
            .O(N__20460),
            .I(\sb_translator_1.cnt_leds_RNITAVEZ0Z_8 ));
    Odrv4 I__4288 (
            .O(N__20457),
            .I(\sb_translator_1.cnt_leds_RNITAVEZ0Z_8 ));
    InMux I__4287 (
            .O(N__20452),
            .I(bfn_8_4_0_));
    InMux I__4286 (
            .O(N__20449),
            .I(N__20446));
    LocalMux I__4285 (
            .O(N__20446),
            .I(N__20443));
    Odrv4 I__4284 (
            .O(N__20443),
            .I(\sb_translator_1.num_leds_RNIH2E91Z0Z_9 ));
    CascadeMux I__4283 (
            .O(N__20440),
            .I(N__20437));
    InMux I__4282 (
            .O(N__20437),
            .I(N__20433));
    InMux I__4281 (
            .O(N__20436),
            .I(N__20430));
    LocalMux I__4280 (
            .O(N__20433),
            .I(N__20427));
    LocalMux I__4279 (
            .O(N__20430),
            .I(\sb_translator_1.num_leds_RNI0EVEZ0Z_8 ));
    Odrv4 I__4278 (
            .O(N__20427),
            .I(\sb_translator_1.num_leds_RNI0EVEZ0Z_8 ));
    InMux I__4277 (
            .O(N__20422),
            .I(\sb_translator_1.state56_a_5_cry_7 ));
    InMux I__4276 (
            .O(N__20419),
            .I(N__20416));
    LocalMux I__4275 (
            .O(N__20416),
            .I(N__20413));
    Odrv4 I__4274 (
            .O(N__20413),
            .I(\sb_translator_1.num_leds_RNICJVN1Z0Z_10 ));
    CascadeMux I__4273 (
            .O(N__20410),
            .I(N__20407));
    InMux I__4272 (
            .O(N__20407),
            .I(N__20404));
    LocalMux I__4271 (
            .O(N__20404),
            .I(N__20401));
    Odrv12 I__4270 (
            .O(N__20401),
            .I(\sb_translator_1.num_leds_RNIHKEQZ0Z_9 ));
    InMux I__4269 (
            .O(N__20398),
            .I(\sb_translator_1.state56_a_5_cry_8 ));
    InMux I__4268 (
            .O(N__20395),
            .I(N__20392));
    LocalMux I__4267 (
            .O(N__20392),
            .I(N__20389));
    Odrv4 I__4266 (
            .O(N__20389),
            .I(\sb_translator_1.num_leds_RNIP02R1Z0Z_11 ));
    CascadeMux I__4265 (
            .O(N__20386),
            .I(N__20383));
    InMux I__4264 (
            .O(N__20383),
            .I(N__20380));
    LocalMux I__4263 (
            .O(N__20380),
            .I(N__20377));
    Odrv12 I__4262 (
            .O(N__20377),
            .I(\sb_translator_1.num_leds_RNIRUGTZ0Z_10 ));
    InMux I__4261 (
            .O(N__20374),
            .I(\sb_translator_1.state56_a_5_cry_9 ));
    InMux I__4260 (
            .O(N__20371),
            .I(\sb_translator_1.state56_a_5_cry_10 ));
    InMux I__4259 (
            .O(N__20368),
            .I(\sb_translator_1.state56_a_5_cry_11 ));
    CascadeMux I__4258 (
            .O(N__20365),
            .I(N__20362));
    InMux I__4257 (
            .O(N__20362),
            .I(N__20355));
    InMux I__4256 (
            .O(N__20361),
            .I(N__20348));
    InMux I__4255 (
            .O(N__20360),
            .I(N__20348));
    InMux I__4254 (
            .O(N__20359),
            .I(N__20348));
    InMux I__4253 (
            .O(N__20358),
            .I(N__20345));
    LocalMux I__4252 (
            .O(N__20355),
            .I(N__20342));
    LocalMux I__4251 (
            .O(N__20348),
            .I(N__20339));
    LocalMux I__4250 (
            .O(N__20345),
            .I(N__20336));
    Span4Mux_v I__4249 (
            .O(N__20342),
            .I(N__20333));
    Span4Mux_v I__4248 (
            .O(N__20339),
            .I(N__20330));
    Span4Mux_h I__4247 (
            .O(N__20336),
            .I(N__20327));
    Odrv4 I__4246 (
            .O(N__20333),
            .I(ram_sel_13));
    Odrv4 I__4245 (
            .O(N__20330),
            .I(ram_sel_13));
    Odrv4 I__4244 (
            .O(N__20327),
            .I(ram_sel_13));
    CascadeMux I__4243 (
            .O(N__20320),
            .I(N__20313));
    InMux I__4242 (
            .O(N__20319),
            .I(N__20309));
    InMux I__4241 (
            .O(N__20318),
            .I(N__20302));
    InMux I__4240 (
            .O(N__20317),
            .I(N__20302));
    InMux I__4239 (
            .O(N__20316),
            .I(N__20302));
    InMux I__4238 (
            .O(N__20313),
            .I(N__20297));
    InMux I__4237 (
            .O(N__20312),
            .I(N__20297));
    LocalMux I__4236 (
            .O(N__20309),
            .I(N__20294));
    LocalMux I__4235 (
            .O(N__20302),
            .I(N__20291));
    LocalMux I__4234 (
            .O(N__20297),
            .I(N__20288));
    Span4Mux_v I__4233 (
            .O(N__20294),
            .I(N__20283));
    Span4Mux_v I__4232 (
            .O(N__20291),
            .I(N__20283));
    Span4Mux_h I__4231 (
            .O(N__20288),
            .I(N__20280));
    Odrv4 I__4230 (
            .O(N__20283),
            .I(ram_sel_10));
    Odrv4 I__4229 (
            .O(N__20280),
            .I(ram_sel_10));
    CascadeMux I__4228 (
            .O(N__20275),
            .I(N__20270));
    InMux I__4227 (
            .O(N__20274),
            .I(N__20264));
    InMux I__4226 (
            .O(N__20273),
            .I(N__20259));
    InMux I__4225 (
            .O(N__20270),
            .I(N__20259));
    InMux I__4224 (
            .O(N__20269),
            .I(N__20254));
    InMux I__4223 (
            .O(N__20268),
            .I(N__20254));
    InMux I__4222 (
            .O(N__20267),
            .I(N__20251));
    LocalMux I__4221 (
            .O(N__20264),
            .I(N__20246));
    LocalMux I__4220 (
            .O(N__20259),
            .I(N__20246));
    LocalMux I__4219 (
            .O(N__20254),
            .I(N__20243));
    LocalMux I__4218 (
            .O(N__20251),
            .I(N__20240));
    Span4Mux_h I__4217 (
            .O(N__20246),
            .I(N__20237));
    Span4Mux_h I__4216 (
            .O(N__20243),
            .I(N__20234));
    Odrv4 I__4215 (
            .O(N__20240),
            .I(ram_sel_7));
    Odrv4 I__4214 (
            .O(N__20237),
            .I(ram_sel_7));
    Odrv4 I__4213 (
            .O(N__20234),
            .I(ram_sel_7));
    CascadeMux I__4212 (
            .O(N__20227),
            .I(N__20223));
    CascadeMux I__4211 (
            .O(N__20226),
            .I(N__20218));
    InMux I__4210 (
            .O(N__20223),
            .I(N__20212));
    InMux I__4209 (
            .O(N__20222),
            .I(N__20212));
    InMux I__4208 (
            .O(N__20221),
            .I(N__20209));
    InMux I__4207 (
            .O(N__20218),
            .I(N__20204));
    InMux I__4206 (
            .O(N__20217),
            .I(N__20204));
    LocalMux I__4205 (
            .O(N__20212),
            .I(\demux.N_240 ));
    LocalMux I__4204 (
            .O(N__20209),
            .I(\demux.N_240 ));
    LocalMux I__4203 (
            .O(N__20204),
            .I(\demux.N_240 ));
    InMux I__4202 (
            .O(N__20197),
            .I(N__20194));
    LocalMux I__4201 (
            .O(N__20194),
            .I(N__20191));
    Span4Mux_v I__4200 (
            .O(N__20191),
            .I(N__20188));
    Span4Mux_h I__4199 (
            .O(N__20188),
            .I(N__20185));
    Span4Mux_v I__4198 (
            .O(N__20185),
            .I(N__20182));
    Odrv4 I__4197 (
            .O(N__20182),
            .I(demux_data_in_29));
    CascadeMux I__4196 (
            .O(N__20179),
            .I(N__20176));
    InMux I__4195 (
            .O(N__20176),
            .I(N__20173));
    LocalMux I__4194 (
            .O(N__20173),
            .I(N__20169));
    InMux I__4193 (
            .O(N__20172),
            .I(N__20166));
    Span4Mux_s2_v I__4192 (
            .O(N__20169),
            .I(N__20161));
    LocalMux I__4191 (
            .O(N__20166),
            .I(N__20161));
    Odrv4 I__4190 (
            .O(N__20161),
            .I(\sb_translator_1.state56_a_5_ac0_1 ));
    InMux I__4189 (
            .O(N__20158),
            .I(N__20155));
    LocalMux I__4188 (
            .O(N__20155),
            .I(\sb_translator_1.cnt_leds_RNIJDTTZ0Z_2 ));
    CascadeMux I__4187 (
            .O(N__20152),
            .I(N__20149));
    InMux I__4186 (
            .O(N__20149),
            .I(N__20146));
    LocalMux I__4185 (
            .O(N__20146),
            .I(\sb_translator_1.state56_a_5_44 ));
    InMux I__4184 (
            .O(N__20143),
            .I(\sb_translator_1.state56_a_5_cry_0_c_THRU_CO ));
    InMux I__4183 (
            .O(N__20140),
            .I(N__20137));
    LocalMux I__4182 (
            .O(N__20137),
            .I(\sb_translator_1.cnt_leds_RNIBOUEZ0Z_2 ));
    CascadeMux I__4181 (
            .O(N__20134),
            .I(N__20131));
    InMux I__4180 (
            .O(N__20131),
            .I(N__20128));
    LocalMux I__4179 (
            .O(N__20128),
            .I(\sb_translator_1.cnt_leds_RNIPJTTZ0Z_3 ));
    InMux I__4178 (
            .O(N__20125),
            .I(\sb_translator_1.state56_a_5_cry_0 ));
    InMux I__4177 (
            .O(N__20122),
            .I(N__20119));
    LocalMux I__4176 (
            .O(N__20119),
            .I(\sb_translator_1.cnt_leds_RNIERUEZ0Z_3 ));
    CascadeMux I__4175 (
            .O(N__20116),
            .I(N__20113));
    InMux I__4174 (
            .O(N__20113),
            .I(N__20110));
    LocalMux I__4173 (
            .O(N__20110),
            .I(\sb_translator_1.cnt_leds_RNIVPTTZ0Z_4 ));
    InMux I__4172 (
            .O(N__20107),
            .I(\sb_translator_1.state56_a_5_cry_1 ));
    InMux I__4171 (
            .O(N__20104),
            .I(N__20100));
    InMux I__4170 (
            .O(N__20103),
            .I(N__20097));
    LocalMux I__4169 (
            .O(N__20100),
            .I(\sb_translator_1.cnt_leds_RNIHUUEZ0Z_4 ));
    LocalMux I__4168 (
            .O(N__20097),
            .I(\sb_translator_1.cnt_leds_RNIHUUEZ0Z_4 ));
    CascadeMux I__4167 (
            .O(N__20092),
            .I(N__20089));
    InMux I__4166 (
            .O(N__20089),
            .I(N__20086));
    LocalMux I__4165 (
            .O(N__20086),
            .I(\sb_translator_1.cnt_leds_RNI50UTZ0Z_5 ));
    InMux I__4164 (
            .O(N__20083),
            .I(\sb_translator_1.state56_a_5_cry_2 ));
    InMux I__4163 (
            .O(N__20080),
            .I(N__20077));
    LocalMux I__4162 (
            .O(N__20077),
            .I(\sb_translator_1.cnt_leds_RNIK1VEZ0Z_5 ));
    CascadeMux I__4161 (
            .O(N__20074),
            .I(N__20071));
    InMux I__4160 (
            .O(N__20071),
            .I(N__20068));
    LocalMux I__4159 (
            .O(N__20068),
            .I(\sb_translator_1.cnt_leds_RNIB6UTZ0Z_6 ));
    InMux I__4158 (
            .O(N__20065),
            .I(\sb_translator_1.state56_a_5_cry_3 ));
    InMux I__4157 (
            .O(N__20062),
            .I(N__20059));
    LocalMux I__4156 (
            .O(N__20059),
            .I(\demux.N_917 ));
    CascadeMux I__4155 (
            .O(N__20056),
            .I(\demux.N_424_i_0_o2_0_7_cascade_ ));
    InMux I__4154 (
            .O(N__20053),
            .I(N__20050));
    LocalMux I__4153 (
            .O(N__20050),
            .I(\demux.N_424_i_0_o2_0_10 ));
    CascadeMux I__4152 (
            .O(N__20047),
            .I(\demux.N_424_i_0_o2Z0Z_0_cascade_ ));
    InMux I__4151 (
            .O(N__20044),
            .I(N__20041));
    LocalMux I__4150 (
            .O(N__20041),
            .I(N__20038));
    Span4Mux_h I__4149 (
            .O(N__20038),
            .I(N__20035));
    Odrv4 I__4148 (
            .O(N__20035),
            .I(demux_data_in_16));
    CascadeMux I__4147 (
            .O(N__20032),
            .I(N__20029));
    InMux I__4146 (
            .O(N__20029),
            .I(N__20026));
    LocalMux I__4145 (
            .O(N__20026),
            .I(N__20023));
    Span4Mux_h I__4144 (
            .O(N__20023),
            .I(N__20020));
    Odrv4 I__4143 (
            .O(N__20020),
            .I(demux_data_in_96));
    InMux I__4142 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__4141 (
            .O(N__20014),
            .I(N__20011));
    Span4Mux_h I__4140 (
            .O(N__20011),
            .I(N__20008));
    Odrv4 I__4139 (
            .O(N__20008),
            .I(demux_data_in_64));
    CascadeMux I__4138 (
            .O(N__20005),
            .I(\demux.N_424_i_0_o2Z0Z_4_cascade_ ));
    InMux I__4137 (
            .O(N__20002),
            .I(N__19998));
    InMux I__4136 (
            .O(N__20001),
            .I(N__19995));
    LocalMux I__4135 (
            .O(N__19998),
            .I(N__19991));
    LocalMux I__4134 (
            .O(N__19995),
            .I(N__19988));
    InMux I__4133 (
            .O(N__19994),
            .I(N__19985));
    Span4Mux_h I__4132 (
            .O(N__19991),
            .I(N__19978));
    Span4Mux_h I__4131 (
            .O(N__19988),
            .I(N__19978));
    LocalMux I__4130 (
            .O(N__19985),
            .I(N__19978));
    Odrv4 I__4129 (
            .O(N__19978),
            .I(\demux.N_424_i_0_o2Z0Z_8 ));
    InMux I__4128 (
            .O(N__19975),
            .I(N__19972));
    LocalMux I__4127 (
            .O(N__19972),
            .I(N__19967));
    InMux I__4126 (
            .O(N__19971),
            .I(N__19964));
    CascadeMux I__4125 (
            .O(N__19970),
            .I(N__19961));
    Span4Mux_v I__4124 (
            .O(N__19967),
            .I(N__19956));
    LocalMux I__4123 (
            .O(N__19964),
            .I(N__19956));
    InMux I__4122 (
            .O(N__19961),
            .I(N__19953));
    Odrv4 I__4121 (
            .O(N__19956),
            .I(\demux.N_424_i_0_aZ0Z3 ));
    LocalMux I__4120 (
            .O(N__19953),
            .I(\demux.N_424_i_0_aZ0Z3 ));
    InMux I__4119 (
            .O(N__19948),
            .I(N__19944));
    InMux I__4118 (
            .O(N__19947),
            .I(N__19941));
    LocalMux I__4117 (
            .O(N__19944),
            .I(N__19937));
    LocalMux I__4116 (
            .O(N__19941),
            .I(N__19934));
    InMux I__4115 (
            .O(N__19940),
            .I(N__19931));
    Span4Mux_h I__4114 (
            .O(N__19937),
            .I(N__19925));
    Span4Mux_h I__4113 (
            .O(N__19934),
            .I(N__19925));
    LocalMux I__4112 (
            .O(N__19931),
            .I(N__19922));
    InMux I__4111 (
            .O(N__19930),
            .I(N__19919));
    Odrv4 I__4110 (
            .O(N__19925),
            .I(\demux.N_424_i_0_o2_9 ));
    Odrv4 I__4109 (
            .O(N__19922),
            .I(\demux.N_424_i_0_o2_9 ));
    LocalMux I__4108 (
            .O(N__19919),
            .I(\demux.N_424_i_0_o2_9 ));
    CascadeMux I__4107 (
            .O(N__19912),
            .I(\demux.N_424_i_0_o2Z0Z_8_cascade_ ));
    InMux I__4106 (
            .O(N__19909),
            .I(N__19905));
    CascadeMux I__4105 (
            .O(N__19908),
            .I(N__19902));
    LocalMux I__4104 (
            .O(N__19905),
            .I(N__19899));
    InMux I__4103 (
            .O(N__19902),
            .I(N__19896));
    Span4Mux_v I__4102 (
            .O(N__19899),
            .I(N__19889));
    LocalMux I__4101 (
            .O(N__19896),
            .I(N__19889));
    InMux I__4100 (
            .O(N__19895),
            .I(N__19886));
    InMux I__4099 (
            .O(N__19894),
            .I(N__19883));
    Odrv4 I__4098 (
            .O(N__19889),
            .I(\demux.N_424_i_0_o2Z0Z_7 ));
    LocalMux I__4097 (
            .O(N__19886),
            .I(\demux.N_424_i_0_o2Z0Z_7 ));
    LocalMux I__4096 (
            .O(N__19883),
            .I(\demux.N_424_i_0_o2Z0Z_7 ));
    InMux I__4095 (
            .O(N__19876),
            .I(N__19873));
    LocalMux I__4094 (
            .O(N__19873),
            .I(N__19870));
    Span4Mux_v I__4093 (
            .O(N__19870),
            .I(N__19867));
    Span4Mux_h I__4092 (
            .O(N__19867),
            .I(N__19864));
    Span4Mux_v I__4091 (
            .O(N__19864),
            .I(N__19861));
    Odrv4 I__4090 (
            .O(N__19861),
            .I(demux_data_in_24));
    InMux I__4089 (
            .O(N__19858),
            .I(N__19855));
    LocalMux I__4088 (
            .O(N__19855),
            .I(\demux.N_424_i_0_a3Z0Z_7 ));
    InMux I__4087 (
            .O(N__19852),
            .I(N__19849));
    LocalMux I__4086 (
            .O(N__19849),
            .I(N__19845));
    CascadeMux I__4085 (
            .O(N__19848),
            .I(N__19841));
    Span4Mux_v I__4084 (
            .O(N__19845),
            .I(N__19837));
    InMux I__4083 (
            .O(N__19844),
            .I(N__19834));
    InMux I__4082 (
            .O(N__19841),
            .I(N__19831));
    InMux I__4081 (
            .O(N__19840),
            .I(N__19828));
    Odrv4 I__4080 (
            .O(N__19837),
            .I(ram_sel_0));
    LocalMux I__4079 (
            .O(N__19834),
            .I(ram_sel_0));
    LocalMux I__4078 (
            .O(N__19831),
            .I(ram_sel_0));
    LocalMux I__4077 (
            .O(N__19828),
            .I(ram_sel_0));
    InMux I__4076 (
            .O(N__19819),
            .I(N__19814));
    CascadeMux I__4075 (
            .O(N__19818),
            .I(N__19811));
    InMux I__4074 (
            .O(N__19817),
            .I(N__19807));
    LocalMux I__4073 (
            .O(N__19814),
            .I(N__19803));
    InMux I__4072 (
            .O(N__19811),
            .I(N__19798));
    InMux I__4071 (
            .O(N__19810),
            .I(N__19798));
    LocalMux I__4070 (
            .O(N__19807),
            .I(N__19795));
    InMux I__4069 (
            .O(N__19806),
            .I(N__19792));
    Span4Mux_v I__4068 (
            .O(N__19803),
            .I(N__19789));
    LocalMux I__4067 (
            .O(N__19798),
            .I(N__19786));
    Span4Mux_h I__4066 (
            .O(N__19795),
            .I(N__19783));
    LocalMux I__4065 (
            .O(N__19792),
            .I(N__19780));
    Odrv4 I__4064 (
            .O(N__19789),
            .I(ram_sel_11));
    Odrv4 I__4063 (
            .O(N__19786),
            .I(ram_sel_11));
    Odrv4 I__4062 (
            .O(N__19783),
            .I(ram_sel_11));
    Odrv12 I__4061 (
            .O(N__19780),
            .I(ram_sel_11));
    CascadeMux I__4060 (
            .O(N__19771),
            .I(\demux.N_906_cascade_ ));
    InMux I__4059 (
            .O(N__19768),
            .I(N__19764));
    InMux I__4058 (
            .O(N__19767),
            .I(N__19761));
    LocalMux I__4057 (
            .O(N__19764),
            .I(N__19758));
    LocalMux I__4056 (
            .O(N__19761),
            .I(N__19753));
    Span4Mux_v I__4055 (
            .O(N__19758),
            .I(N__19749));
    InMux I__4054 (
            .O(N__19757),
            .I(N__19744));
    InMux I__4053 (
            .O(N__19756),
            .I(N__19744));
    Span4Mux_h I__4052 (
            .O(N__19753),
            .I(N__19741));
    InMux I__4051 (
            .O(N__19752),
            .I(N__19738));
    Odrv4 I__4050 (
            .O(N__19749),
            .I(ram_sel_4));
    LocalMux I__4049 (
            .O(N__19744),
            .I(ram_sel_4));
    Odrv4 I__4048 (
            .O(N__19741),
            .I(ram_sel_4));
    LocalMux I__4047 (
            .O(N__19738),
            .I(ram_sel_4));
    InMux I__4046 (
            .O(N__19729),
            .I(N__19726));
    LocalMux I__4045 (
            .O(N__19726),
            .I(\demux.N_424_i_0_o2_0Z0Z_3 ));
    InMux I__4044 (
            .O(N__19723),
            .I(N__19720));
    LocalMux I__4043 (
            .O(N__19720),
            .I(N__19717));
    Span4Mux_v I__4042 (
            .O(N__19717),
            .I(N__19714));
    Span4Mux_h I__4041 (
            .O(N__19714),
            .I(N__19711));
    Span4Mux_v I__4040 (
            .O(N__19711),
            .I(N__19708));
    Odrv4 I__4039 (
            .O(N__19708),
            .I(demux_data_in_28));
    CascadeMux I__4038 (
            .O(N__19705),
            .I(\demux.N_918_cascade_ ));
    InMux I__4037 (
            .O(N__19702),
            .I(N__19699));
    LocalMux I__4036 (
            .O(N__19699),
            .I(N__19696));
    Span4Mux_h I__4035 (
            .O(N__19696),
            .I(N__19693));
    Odrv4 I__4034 (
            .O(N__19693),
            .I(demux_data_in_105));
    CascadeMux I__4033 (
            .O(N__19690),
            .I(\demux.N_424_i_0_a2Z0Z_5_cascade_ ));
    InMux I__4032 (
            .O(N__19687),
            .I(N__19684));
    LocalMux I__4031 (
            .O(N__19684),
            .I(N__19681));
    Span4Mux_v I__4030 (
            .O(N__19681),
            .I(N__19678));
    Span4Mux_h I__4029 (
            .O(N__19678),
            .I(N__19675));
    Odrv4 I__4028 (
            .O(N__19675),
            .I(demux_data_in_33));
    InMux I__4027 (
            .O(N__19672),
            .I(N__19669));
    LocalMux I__4026 (
            .O(N__19669),
            .I(\demux.N_423_i_0_o2Z0Z_0 ));
    InMux I__4025 (
            .O(N__19666),
            .I(N__19662));
    InMux I__4024 (
            .O(N__19665),
            .I(N__19659));
    LocalMux I__4023 (
            .O(N__19662),
            .I(\demux.N_918 ));
    LocalMux I__4022 (
            .O(N__19659),
            .I(\demux.N_918 ));
    InMux I__4021 (
            .O(N__19654),
            .I(N__19646));
    InMux I__4020 (
            .O(N__19653),
            .I(N__19646));
    InMux I__4019 (
            .O(N__19652),
            .I(N__19637));
    InMux I__4018 (
            .O(N__19651),
            .I(N__19637));
    LocalMux I__4017 (
            .O(N__19646),
            .I(N__19634));
    InMux I__4016 (
            .O(N__19645),
            .I(N__19625));
    InMux I__4015 (
            .O(N__19644),
            .I(N__19625));
    InMux I__4014 (
            .O(N__19643),
            .I(N__19625));
    InMux I__4013 (
            .O(N__19642),
            .I(N__19625));
    LocalMux I__4012 (
            .O(N__19637),
            .I(N__19618));
    Span4Mux_v I__4011 (
            .O(N__19634),
            .I(N__19618));
    LocalMux I__4010 (
            .O(N__19625),
            .I(N__19618));
    Odrv4 I__4009 (
            .O(N__19618),
            .I(\demux.N_424_i_0_a2Z0Z_7 ));
    InMux I__4008 (
            .O(N__19615),
            .I(N__19612));
    LocalMux I__4007 (
            .O(N__19612),
            .I(N__19609));
    Span4Mux_h I__4006 (
            .O(N__19609),
            .I(N__19606));
    Odrv4 I__4005 (
            .O(N__19606),
            .I(\demux.N_424_i_0_o2_0_1 ));
    InMux I__4004 (
            .O(N__19603),
            .I(N__19599));
    CascadeMux I__4003 (
            .O(N__19602),
            .I(N__19596));
    LocalMux I__4002 (
            .O(N__19599),
            .I(N__19592));
    InMux I__4001 (
            .O(N__19596),
            .I(N__19587));
    InMux I__4000 (
            .O(N__19595),
            .I(N__19587));
    Span4Mux_v I__3999 (
            .O(N__19592),
            .I(N__19584));
    LocalMux I__3998 (
            .O(N__19587),
            .I(N__19579));
    Span4Mux_h I__3997 (
            .O(N__19584),
            .I(N__19579));
    Odrv4 I__3996 (
            .O(N__19579),
            .I(\demux.N_236 ));
    InMux I__3995 (
            .O(N__19576),
            .I(N__19573));
    LocalMux I__3994 (
            .O(N__19573),
            .I(N__19570));
    Span4Mux_h I__3993 (
            .O(N__19570),
            .I(N__19566));
    InMux I__3992 (
            .O(N__19569),
            .I(N__19563));
    Odrv4 I__3991 (
            .O(N__19566),
            .I(\demux.N_235 ));
    LocalMux I__3990 (
            .O(N__19563),
            .I(\demux.N_235 ));
    InMux I__3989 (
            .O(N__19558),
            .I(N__19555));
    LocalMux I__3988 (
            .O(N__19555),
            .I(\demux.N_424_i_0_o2_0Z0Z_2 ));
    InMux I__3987 (
            .O(N__19552),
            .I(N__19547));
    InMux I__3986 (
            .O(N__19551),
            .I(N__19542));
    InMux I__3985 (
            .O(N__19550),
            .I(N__19542));
    LocalMux I__3984 (
            .O(N__19547),
            .I(\demux.N_237 ));
    LocalMux I__3983 (
            .O(N__19542),
            .I(\demux.N_237 ));
    CascadeMux I__3982 (
            .O(N__19537),
            .I(\demux.N_424_i_0_o2_0_8Z0Z_1_cascade_ ));
    InMux I__3981 (
            .O(N__19534),
            .I(N__19529));
    InMux I__3980 (
            .O(N__19533),
            .I(N__19524));
    InMux I__3979 (
            .O(N__19532),
            .I(N__19524));
    LocalMux I__3978 (
            .O(N__19529),
            .I(\demux.N_238 ));
    LocalMux I__3977 (
            .O(N__19524),
            .I(\demux.N_238 ));
    InMux I__3976 (
            .O(N__19519),
            .I(N__19516));
    LocalMux I__3975 (
            .O(N__19516),
            .I(N__19513));
    Span4Mux_v I__3974 (
            .O(N__19513),
            .I(N__19510));
    Odrv4 I__3973 (
            .O(N__19510),
            .I(demux_data_in_91));
    CascadeMux I__3972 (
            .O(N__19507),
            .I(\demux.N_421_i_0_o2Z0Z_0_cascade_ ));
    InMux I__3971 (
            .O(N__19504),
            .I(N__19501));
    LocalMux I__3970 (
            .O(N__19501),
            .I(N__19498));
    Span4Mux_v I__3969 (
            .O(N__19498),
            .I(N__19495));
    Span4Mux_h I__3968 (
            .O(N__19495),
            .I(N__19492));
    Odrv4 I__3967 (
            .O(N__19492),
            .I(demux_data_in_2));
    InMux I__3966 (
            .O(N__19489),
            .I(N__19486));
    LocalMux I__3965 (
            .O(N__19486),
            .I(N__19483));
    Span4Mux_v I__3964 (
            .O(N__19483),
            .I(N__19480));
    Odrv4 I__3963 (
            .O(N__19480),
            .I(demux_data_in_106));
    InMux I__3962 (
            .O(N__19477),
            .I(N__19474));
    LocalMux I__3961 (
            .O(N__19474),
            .I(N__19471));
    Span4Mux_v I__3960 (
            .O(N__19471),
            .I(N__19468));
    Odrv4 I__3959 (
            .O(N__19468),
            .I(demux_data_in_34));
    CascadeMux I__3958 (
            .O(N__19465),
            .I(\demux.N_422_i_0_o2Z0Z_0_cascade_ ));
    InMux I__3957 (
            .O(N__19462),
            .I(N__19459));
    LocalMux I__3956 (
            .O(N__19459),
            .I(N__19456));
    Span4Mux_v I__3955 (
            .O(N__19456),
            .I(N__19453));
    Odrv4 I__3954 (
            .O(N__19453),
            .I(demux_data_in_90));
    InMux I__3953 (
            .O(N__19450),
            .I(N__19447));
    LocalMux I__3952 (
            .O(N__19447),
            .I(\demux.N_422_i_0_a3Z0Z_4 ));
    InMux I__3951 (
            .O(N__19444),
            .I(N__19441));
    LocalMux I__3950 (
            .O(N__19441),
            .I(N__19438));
    Span4Mux_h I__3949 (
            .O(N__19438),
            .I(N__19435));
    Odrv4 I__3948 (
            .O(N__19435),
            .I(demux_data_in_10));
    CascadeMux I__3947 (
            .O(N__19432),
            .I(\demux.N_422_i_0_o2Z0Z_1_cascade_ ));
    InMux I__3946 (
            .O(N__19429),
            .I(N__19426));
    LocalMux I__3945 (
            .O(N__19426),
            .I(N__19423));
    Span4Mux_v I__3944 (
            .O(N__19423),
            .I(N__19420));
    Odrv4 I__3943 (
            .O(N__19420),
            .I(demux_data_in_9));
    InMux I__3942 (
            .O(N__19417),
            .I(N__19414));
    LocalMux I__3941 (
            .O(N__19414),
            .I(N__19411));
    Span4Mux_v I__3940 (
            .O(N__19411),
            .I(N__19408));
    Odrv4 I__3939 (
            .O(N__19408),
            .I(demux_data_in_89));
    CascadeMux I__3938 (
            .O(N__19405),
            .I(\demux.N_423_i_0_a3Z0Z_5_cascade_ ));
    InMux I__3937 (
            .O(N__19402),
            .I(N__19399));
    LocalMux I__3936 (
            .O(N__19399),
            .I(N__19396));
    Span4Mux_v I__3935 (
            .O(N__19396),
            .I(N__19393));
    Odrv4 I__3934 (
            .O(N__19393),
            .I(demux_data_in_43));
    InMux I__3933 (
            .O(N__19390),
            .I(N__19387));
    LocalMux I__3932 (
            .O(N__19387),
            .I(\demux.N_837 ));
    InMux I__3931 (
            .O(N__19384),
            .I(N__19380));
    InMux I__3930 (
            .O(N__19383),
            .I(N__19377));
    LocalMux I__3929 (
            .O(N__19380),
            .I(\demux.N_424_i_0_a2Z0Z_34 ));
    LocalMux I__3928 (
            .O(N__19377),
            .I(\demux.N_424_i_0_a2Z0Z_34 ));
    InMux I__3927 (
            .O(N__19372),
            .I(\sb_translator_1.cnt_leds_cry_14 ));
    InMux I__3926 (
            .O(N__19369),
            .I(bfn_7_6_0_));
    CEMux I__3925 (
            .O(N__19366),
            .I(N__19362));
    CEMux I__3924 (
            .O(N__19365),
            .I(N__19359));
    LocalMux I__3923 (
            .O(N__19362),
            .I(N__19356));
    LocalMux I__3922 (
            .O(N__19359),
            .I(N__19352));
    Span4Mux_v I__3921 (
            .O(N__19356),
            .I(N__19349));
    CEMux I__3920 (
            .O(N__19355),
            .I(N__19346));
    Odrv4 I__3919 (
            .O(N__19352),
            .I(\sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1 ));
    Odrv4 I__3918 (
            .O(N__19349),
            .I(\sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1 ));
    LocalMux I__3917 (
            .O(N__19346),
            .I(\sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1 ));
    InMux I__3916 (
            .O(N__19339),
            .I(N__19336));
    LocalMux I__3915 (
            .O(N__19336),
            .I(N__19333));
    Span4Mux_h I__3914 (
            .O(N__19333),
            .I(N__19330));
    Odrv4 I__3913 (
            .O(N__19330),
            .I(demux_data_in_40));
    InMux I__3912 (
            .O(N__19327),
            .I(N__19324));
    LocalMux I__3911 (
            .O(N__19324),
            .I(N__19321));
    Span4Mux_v I__3910 (
            .O(N__19321),
            .I(N__19318));
    Odrv4 I__3909 (
            .O(N__19318),
            .I(demux_data_in_88));
    InMux I__3908 (
            .O(N__19315),
            .I(N__19312));
    LocalMux I__3907 (
            .O(N__19312),
            .I(\demux.N_424_i_0_a3Z0Z_4 ));
    InMux I__3906 (
            .O(N__19309),
            .I(N__19306));
    LocalMux I__3905 (
            .O(N__19306),
            .I(N__19303));
    Span4Mux_h I__3904 (
            .O(N__19303),
            .I(N__19300));
    Span4Mux_v I__3903 (
            .O(N__19300),
            .I(N__19297));
    Odrv4 I__3902 (
            .O(N__19297),
            .I(demux_data_in_8));
    CascadeMux I__3901 (
            .O(N__19294),
            .I(\demux.N_424_i_0_o2Z0Z_1_cascade_ ));
    InMux I__3900 (
            .O(N__19291),
            .I(N__19288));
    LocalMux I__3899 (
            .O(N__19288),
            .I(N__19285));
    Span4Mux_h I__3898 (
            .O(N__19285),
            .I(N__19282));
    Span4Mux_v I__3897 (
            .O(N__19282),
            .I(N__19279));
    Odrv4 I__3896 (
            .O(N__19279),
            .I(demux_data_in_0));
    CascadeMux I__3895 (
            .O(N__19276),
            .I(\demux.N_424_i_0_aZ0Z3_cascade_ ));
    InMux I__3894 (
            .O(N__19273),
            .I(N__19270));
    LocalMux I__3893 (
            .O(N__19270),
            .I(N__19267));
    Span4Mux_v I__3892 (
            .O(N__19267),
            .I(N__19264));
    Odrv4 I__3891 (
            .O(N__19264),
            .I(demux_data_in_35));
    CascadeMux I__3890 (
            .O(N__19261),
            .I(N__19258));
    InMux I__3889 (
            .O(N__19258),
            .I(N__19255));
    LocalMux I__3888 (
            .O(N__19255),
            .I(N__19252));
    Span4Mux_h I__3887 (
            .O(N__19252),
            .I(N__19249));
    Odrv4 I__3886 (
            .O(N__19249),
            .I(demux_data_in_107));
    InMux I__3885 (
            .O(N__19246),
            .I(N__19238));
    InMux I__3884 (
            .O(N__19245),
            .I(N__19238));
    InMux I__3883 (
            .O(N__19244),
            .I(N__19235));
    InMux I__3882 (
            .O(N__19243),
            .I(N__19232));
    LocalMux I__3881 (
            .O(N__19238),
            .I(N__19229));
    LocalMux I__3880 (
            .O(N__19235),
            .I(\sb_translator_1.cnt_ledsZ0Z_7 ));
    LocalMux I__3879 (
            .O(N__19232),
            .I(\sb_translator_1.cnt_ledsZ0Z_7 ));
    Odrv4 I__3878 (
            .O(N__19229),
            .I(\sb_translator_1.cnt_ledsZ0Z_7 ));
    InMux I__3877 (
            .O(N__19222),
            .I(\sb_translator_1.cnt_leds_cry_6 ));
    InMux I__3876 (
            .O(N__19219),
            .I(N__19216));
    LocalMux I__3875 (
            .O(N__19216),
            .I(N__19210));
    InMux I__3874 (
            .O(N__19215),
            .I(N__19205));
    InMux I__3873 (
            .O(N__19214),
            .I(N__19205));
    InMux I__3872 (
            .O(N__19213),
            .I(N__19202));
    Sp12to4 I__3871 (
            .O(N__19210),
            .I(N__19197));
    LocalMux I__3870 (
            .O(N__19205),
            .I(N__19197));
    LocalMux I__3869 (
            .O(N__19202),
            .I(\sb_translator_1.cnt_ledsZ0Z_8 ));
    Odrv12 I__3868 (
            .O(N__19197),
            .I(\sb_translator_1.cnt_ledsZ0Z_8 ));
    InMux I__3867 (
            .O(N__19192),
            .I(bfn_7_5_0_));
    InMux I__3866 (
            .O(N__19189),
            .I(\sb_translator_1.cnt_leds_cry_8 ));
    InMux I__3865 (
            .O(N__19186),
            .I(N__19177));
    InMux I__3864 (
            .O(N__19185),
            .I(N__19172));
    InMux I__3863 (
            .O(N__19184),
            .I(N__19172));
    InMux I__3862 (
            .O(N__19183),
            .I(N__19163));
    InMux I__3861 (
            .O(N__19182),
            .I(N__19163));
    InMux I__3860 (
            .O(N__19181),
            .I(N__19163));
    InMux I__3859 (
            .O(N__19180),
            .I(N__19163));
    LocalMux I__3858 (
            .O(N__19177),
            .I(\sb_translator_1.cnt_ledsZ0Z_10 ));
    LocalMux I__3857 (
            .O(N__19172),
            .I(\sb_translator_1.cnt_ledsZ0Z_10 ));
    LocalMux I__3856 (
            .O(N__19163),
            .I(\sb_translator_1.cnt_ledsZ0Z_10 ));
    InMux I__3855 (
            .O(N__19156),
            .I(\sb_translator_1.cnt_leds_cry_9 ));
    InMux I__3854 (
            .O(N__19153),
            .I(N__19144));
    InMux I__3853 (
            .O(N__19152),
            .I(N__19141));
    InMux I__3852 (
            .O(N__19151),
            .I(N__19138));
    InMux I__3851 (
            .O(N__19150),
            .I(N__19129));
    InMux I__3850 (
            .O(N__19149),
            .I(N__19129));
    InMux I__3849 (
            .O(N__19148),
            .I(N__19129));
    InMux I__3848 (
            .O(N__19147),
            .I(N__19129));
    LocalMux I__3847 (
            .O(N__19144),
            .I(\sb_translator_1.cnt_ledsZ0Z_11 ));
    LocalMux I__3846 (
            .O(N__19141),
            .I(\sb_translator_1.cnt_ledsZ0Z_11 ));
    LocalMux I__3845 (
            .O(N__19138),
            .I(\sb_translator_1.cnt_ledsZ0Z_11 ));
    LocalMux I__3844 (
            .O(N__19129),
            .I(\sb_translator_1.cnt_ledsZ0Z_11 ));
    InMux I__3843 (
            .O(N__19120),
            .I(\sb_translator_1.cnt_leds_cry_10 ));
    InMux I__3842 (
            .O(N__19117),
            .I(\sb_translator_1.cnt_leds_cry_11 ));
    InMux I__3841 (
            .O(N__19114),
            .I(\sb_translator_1.cnt_leds_cry_12 ));
    InMux I__3840 (
            .O(N__19111),
            .I(\sb_translator_1.cnt_leds_cry_13 ));
    InMux I__3839 (
            .O(N__19108),
            .I(N__19105));
    LocalMux I__3838 (
            .O(N__19105),
            .I(N__19101));
    InMux I__3837 (
            .O(N__19104),
            .I(N__19098));
    Span4Mux_h I__3836 (
            .O(N__19101),
            .I(N__19090));
    LocalMux I__3835 (
            .O(N__19098),
            .I(N__19090));
    InMux I__3834 (
            .O(N__19097),
            .I(N__19085));
    InMux I__3833 (
            .O(N__19096),
            .I(N__19085));
    InMux I__3832 (
            .O(N__19095),
            .I(N__19082));
    Odrv4 I__3831 (
            .O(N__19090),
            .I(\sb_translator_1.cnt19 ));
    LocalMux I__3830 (
            .O(N__19085),
            .I(\sb_translator_1.cnt19 ));
    LocalMux I__3829 (
            .O(N__19082),
            .I(\sb_translator_1.cnt19 ));
    InMux I__3828 (
            .O(N__19075),
            .I(N__19062));
    InMux I__3827 (
            .O(N__19074),
            .I(N__19062));
    InMux I__3826 (
            .O(N__19073),
            .I(N__19062));
    InMux I__3825 (
            .O(N__19072),
            .I(N__19062));
    CascadeMux I__3824 (
            .O(N__19071),
            .I(N__19058));
    LocalMux I__3823 (
            .O(N__19062),
            .I(N__19055));
    InMux I__3822 (
            .O(N__19061),
            .I(N__19050));
    InMux I__3821 (
            .O(N__19058),
            .I(N__19050));
    Odrv4 I__3820 (
            .O(N__19055),
            .I(\sb_translator_1.num_ledsZ0Z_2 ));
    LocalMux I__3819 (
            .O(N__19050),
            .I(\sb_translator_1.num_ledsZ0Z_2 ));
    CascadeMux I__3818 (
            .O(N__19045),
            .I(\sb_translator_1.state56_a_5_44_cascade_ ));
    CascadeMux I__3817 (
            .O(N__19042),
            .I(N__19038));
    InMux I__3816 (
            .O(N__19041),
            .I(N__19030));
    InMux I__3815 (
            .O(N__19038),
            .I(N__19030));
    CascadeMux I__3814 (
            .O(N__19037),
            .I(N__19027));
    CascadeMux I__3813 (
            .O(N__19036),
            .I(N__19024));
    CascadeMux I__3812 (
            .O(N__19035),
            .I(N__19020));
    LocalMux I__3811 (
            .O(N__19030),
            .I(N__19016));
    InMux I__3810 (
            .O(N__19027),
            .I(N__19013));
    InMux I__3809 (
            .O(N__19024),
            .I(N__19004));
    InMux I__3808 (
            .O(N__19023),
            .I(N__19004));
    InMux I__3807 (
            .O(N__19020),
            .I(N__19004));
    InMux I__3806 (
            .O(N__19019),
            .I(N__19004));
    Odrv4 I__3805 (
            .O(N__19016),
            .I(\sb_translator_1.num_ledsZ0Z_1 ));
    LocalMux I__3804 (
            .O(N__19013),
            .I(\sb_translator_1.num_ledsZ0Z_1 ));
    LocalMux I__3803 (
            .O(N__19004),
            .I(\sb_translator_1.num_ledsZ0Z_1 ));
    InMux I__3802 (
            .O(N__18997),
            .I(N__18991));
    InMux I__3801 (
            .O(N__18996),
            .I(N__18988));
    InMux I__3800 (
            .O(N__18995),
            .I(N__18985));
    InMux I__3799 (
            .O(N__18994),
            .I(N__18982));
    LocalMux I__3798 (
            .O(N__18991),
            .I(\sb_translator_1.cnt_ledsZ0Z_0 ));
    LocalMux I__3797 (
            .O(N__18988),
            .I(\sb_translator_1.cnt_ledsZ0Z_0 ));
    LocalMux I__3796 (
            .O(N__18985),
            .I(\sb_translator_1.cnt_ledsZ0Z_0 ));
    LocalMux I__3795 (
            .O(N__18982),
            .I(\sb_translator_1.cnt_ledsZ0Z_0 ));
    InMux I__3794 (
            .O(N__18973),
            .I(bfn_7_4_0_));
    InMux I__3793 (
            .O(N__18970),
            .I(N__18963));
    InMux I__3792 (
            .O(N__18969),
            .I(N__18960));
    InMux I__3791 (
            .O(N__18968),
            .I(N__18955));
    InMux I__3790 (
            .O(N__18967),
            .I(N__18955));
    InMux I__3789 (
            .O(N__18966),
            .I(N__18952));
    LocalMux I__3788 (
            .O(N__18963),
            .I(\sb_translator_1.cnt_ledsZ0Z_1 ));
    LocalMux I__3787 (
            .O(N__18960),
            .I(\sb_translator_1.cnt_ledsZ0Z_1 ));
    LocalMux I__3786 (
            .O(N__18955),
            .I(\sb_translator_1.cnt_ledsZ0Z_1 ));
    LocalMux I__3785 (
            .O(N__18952),
            .I(\sb_translator_1.cnt_ledsZ0Z_1 ));
    InMux I__3784 (
            .O(N__18943),
            .I(\sb_translator_1.cnt_leds_cry_0 ));
    InMux I__3783 (
            .O(N__18940),
            .I(N__18934));
    InMux I__3782 (
            .O(N__18939),
            .I(N__18931));
    InMux I__3781 (
            .O(N__18938),
            .I(N__18926));
    InMux I__3780 (
            .O(N__18937),
            .I(N__18926));
    LocalMux I__3779 (
            .O(N__18934),
            .I(\sb_translator_1.cnt_ledsZ0Z_2 ));
    LocalMux I__3778 (
            .O(N__18931),
            .I(\sb_translator_1.cnt_ledsZ0Z_2 ));
    LocalMux I__3777 (
            .O(N__18926),
            .I(\sb_translator_1.cnt_ledsZ0Z_2 ));
    InMux I__3776 (
            .O(N__18919),
            .I(\sb_translator_1.cnt_leds_cry_1 ));
    CascadeMux I__3775 (
            .O(N__18916),
            .I(N__18911));
    InMux I__3774 (
            .O(N__18915),
            .I(N__18907));
    InMux I__3773 (
            .O(N__18914),
            .I(N__18904));
    InMux I__3772 (
            .O(N__18911),
            .I(N__18899));
    InMux I__3771 (
            .O(N__18910),
            .I(N__18899));
    LocalMux I__3770 (
            .O(N__18907),
            .I(\sb_translator_1.cnt_ledsZ0Z_3 ));
    LocalMux I__3769 (
            .O(N__18904),
            .I(\sb_translator_1.cnt_ledsZ0Z_3 ));
    LocalMux I__3768 (
            .O(N__18899),
            .I(\sb_translator_1.cnt_ledsZ0Z_3 ));
    InMux I__3767 (
            .O(N__18892),
            .I(\sb_translator_1.cnt_leds_cry_2 ));
    CascadeMux I__3766 (
            .O(N__18889),
            .I(N__18884));
    InMux I__3765 (
            .O(N__18888),
            .I(N__18880));
    InMux I__3764 (
            .O(N__18887),
            .I(N__18877));
    InMux I__3763 (
            .O(N__18884),
            .I(N__18872));
    InMux I__3762 (
            .O(N__18883),
            .I(N__18872));
    LocalMux I__3761 (
            .O(N__18880),
            .I(\sb_translator_1.cnt_ledsZ0Z_4 ));
    LocalMux I__3760 (
            .O(N__18877),
            .I(\sb_translator_1.cnt_ledsZ0Z_4 ));
    LocalMux I__3759 (
            .O(N__18872),
            .I(\sb_translator_1.cnt_ledsZ0Z_4 ));
    InMux I__3758 (
            .O(N__18865),
            .I(\sb_translator_1.cnt_leds_cry_3 ));
    CascadeMux I__3757 (
            .O(N__18862),
            .I(N__18859));
    InMux I__3756 (
            .O(N__18859),
            .I(N__18851));
    InMux I__3755 (
            .O(N__18858),
            .I(N__18851));
    InMux I__3754 (
            .O(N__18857),
            .I(N__18848));
    InMux I__3753 (
            .O(N__18856),
            .I(N__18845));
    LocalMux I__3752 (
            .O(N__18851),
            .I(N__18842));
    LocalMux I__3751 (
            .O(N__18848),
            .I(\sb_translator_1.cnt_ledsZ0Z_5 ));
    LocalMux I__3750 (
            .O(N__18845),
            .I(\sb_translator_1.cnt_ledsZ0Z_5 ));
    Odrv4 I__3749 (
            .O(N__18842),
            .I(\sb_translator_1.cnt_ledsZ0Z_5 ));
    InMux I__3748 (
            .O(N__18835),
            .I(\sb_translator_1.cnt_leds_cry_4 ));
    InMux I__3747 (
            .O(N__18832),
            .I(N__18824));
    InMux I__3746 (
            .O(N__18831),
            .I(N__18824));
    InMux I__3745 (
            .O(N__18830),
            .I(N__18821));
    InMux I__3744 (
            .O(N__18829),
            .I(N__18818));
    LocalMux I__3743 (
            .O(N__18824),
            .I(N__18815));
    LocalMux I__3742 (
            .O(N__18821),
            .I(\sb_translator_1.cnt_ledsZ0Z_6 ));
    LocalMux I__3741 (
            .O(N__18818),
            .I(\sb_translator_1.cnt_ledsZ0Z_6 ));
    Odrv4 I__3740 (
            .O(N__18815),
            .I(\sb_translator_1.cnt_ledsZ0Z_6 ));
    InMux I__3739 (
            .O(N__18808),
            .I(\sb_translator_1.cnt_leds_cry_5 ));
    CascadeMux I__3738 (
            .O(N__18805),
            .I(N__18801));
    CascadeMux I__3737 (
            .O(N__18804),
            .I(N__18797));
    InMux I__3736 (
            .O(N__18801),
            .I(N__18786));
    InMux I__3735 (
            .O(N__18800),
            .I(N__18786));
    InMux I__3734 (
            .O(N__18797),
            .I(N__18786));
    InMux I__3733 (
            .O(N__18796),
            .I(N__18786));
    CascadeMux I__3732 (
            .O(N__18795),
            .I(N__18782));
    LocalMux I__3731 (
            .O(N__18786),
            .I(N__18779));
    InMux I__3730 (
            .O(N__18785),
            .I(N__18774));
    InMux I__3729 (
            .O(N__18782),
            .I(N__18774));
    Odrv4 I__3728 (
            .O(N__18779),
            .I(\sb_translator_1.num_ledsZ0Z_6 ));
    LocalMux I__3727 (
            .O(N__18774),
            .I(\sb_translator_1.num_ledsZ0Z_6 ));
    CascadeMux I__3726 (
            .O(N__18769),
            .I(\sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_ ));
    InMux I__3725 (
            .O(N__18766),
            .I(N__18754));
    InMux I__3724 (
            .O(N__18765),
            .I(N__18754));
    InMux I__3723 (
            .O(N__18764),
            .I(N__18754));
    InMux I__3722 (
            .O(N__18763),
            .I(N__18754));
    LocalMux I__3721 (
            .O(N__18754),
            .I(N__18750));
    CascadeMux I__3720 (
            .O(N__18753),
            .I(N__18746));
    Span4Mux_s2_v I__3719 (
            .O(N__18750),
            .I(N__18743));
    InMux I__3718 (
            .O(N__18749),
            .I(N__18738));
    InMux I__3717 (
            .O(N__18746),
            .I(N__18738));
    Odrv4 I__3716 (
            .O(N__18743),
            .I(\sb_translator_1.num_ledsZ0Z_7 ));
    LocalMux I__3715 (
            .O(N__18738),
            .I(\sb_translator_1.num_ledsZ0Z_7 ));
    CascadeMux I__3714 (
            .O(N__18733),
            .I(N__18730));
    InMux I__3713 (
            .O(N__18730),
            .I(N__18723));
    InMux I__3712 (
            .O(N__18729),
            .I(N__18723));
    CascadeMux I__3711 (
            .O(N__18728),
            .I(N__18719));
    LocalMux I__3710 (
            .O(N__18723),
            .I(N__18714));
    InMux I__3709 (
            .O(N__18722),
            .I(N__18711));
    InMux I__3708 (
            .O(N__18719),
            .I(N__18708));
    InMux I__3707 (
            .O(N__18718),
            .I(N__18703));
    InMux I__3706 (
            .O(N__18717),
            .I(N__18703));
    Span4Mux_s3_v I__3705 (
            .O(N__18714),
            .I(N__18700));
    LocalMux I__3704 (
            .O(N__18711),
            .I(\sb_translator_1.num_ledsZ0Z_8 ));
    LocalMux I__3703 (
            .O(N__18708),
            .I(\sb_translator_1.num_ledsZ0Z_8 ));
    LocalMux I__3702 (
            .O(N__18703),
            .I(\sb_translator_1.num_ledsZ0Z_8 ));
    Odrv4 I__3701 (
            .O(N__18700),
            .I(\sb_translator_1.num_ledsZ0Z_8 ));
    CascadeMux I__3700 (
            .O(N__18691),
            .I(\sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_ ));
    CascadeMux I__3699 (
            .O(N__18688),
            .I(\sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_ ));
    CascadeMux I__3698 (
            .O(N__18685),
            .I(N__18677));
    InMux I__3697 (
            .O(N__18684),
            .I(N__18668));
    InMux I__3696 (
            .O(N__18683),
            .I(N__18668));
    InMux I__3695 (
            .O(N__18682),
            .I(N__18668));
    InMux I__3694 (
            .O(N__18681),
            .I(N__18668));
    InMux I__3693 (
            .O(N__18680),
            .I(N__18663));
    InMux I__3692 (
            .O(N__18677),
            .I(N__18663));
    LocalMux I__3691 (
            .O(N__18668),
            .I(N__18660));
    LocalMux I__3690 (
            .O(N__18663),
            .I(\sb_translator_1.num_ledsZ0Z_3 ));
    Odrv4 I__3689 (
            .O(N__18660),
            .I(\sb_translator_1.num_ledsZ0Z_3 ));
    CascadeMux I__3688 (
            .O(N__18655),
            .I(N__18652));
    InMux I__3687 (
            .O(N__18652),
            .I(N__18644));
    InMux I__3686 (
            .O(N__18651),
            .I(N__18644));
    InMux I__3685 (
            .O(N__18650),
            .I(N__18638));
    InMux I__3684 (
            .O(N__18649),
            .I(N__18638));
    LocalMux I__3683 (
            .O(N__18644),
            .I(N__18635));
    CascadeMux I__3682 (
            .O(N__18643),
            .I(N__18631));
    LocalMux I__3681 (
            .O(N__18638),
            .I(N__18626));
    Span4Mux_s2_v I__3680 (
            .O(N__18635),
            .I(N__18626));
    InMux I__3679 (
            .O(N__18634),
            .I(N__18621));
    InMux I__3678 (
            .O(N__18631),
            .I(N__18621));
    Odrv4 I__3677 (
            .O(N__18626),
            .I(\sb_translator_1.num_ledsZ0Z_4 ));
    LocalMux I__3676 (
            .O(N__18621),
            .I(\sb_translator_1.num_ledsZ0Z_4 ));
    InMux I__3675 (
            .O(N__18616),
            .I(N__18613));
    LocalMux I__3674 (
            .O(N__18613),
            .I(\spi_slave_1.miso_data_outZ0Z_12 ));
    InMux I__3673 (
            .O(N__18610),
            .I(N__18607));
    LocalMux I__3672 (
            .O(N__18607),
            .I(\spi_slave_1.miso_data_outZ0Z_11 ));
    InMux I__3671 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__3670 (
            .O(N__18601),
            .I(N__18598));
    Odrv4 I__3669 (
            .O(N__18598),
            .I(\spi_slave_1.miso_RNOZ0Z_6 ));
    InMux I__3668 (
            .O(N__18595),
            .I(N__18592));
    LocalMux I__3667 (
            .O(N__18592),
            .I(\spi_slave_1.miso_data_outZ0Z_16 ));
    InMux I__3666 (
            .O(N__18589),
            .I(N__18586));
    LocalMux I__3665 (
            .O(N__18586),
            .I(\spi_slave_1.miso_data_outZ0Z_0 ));
    InMux I__3664 (
            .O(N__18583),
            .I(N__18575));
    InMux I__3663 (
            .O(N__18582),
            .I(N__18575));
    InMux I__3662 (
            .O(N__18581),
            .I(N__18572));
    CascadeMux I__3661 (
            .O(N__18580),
            .I(N__18568));
    LocalMux I__3660 (
            .O(N__18575),
            .I(N__18565));
    LocalMux I__3659 (
            .O(N__18572),
            .I(N__18560));
    InMux I__3658 (
            .O(N__18571),
            .I(N__18557));
    InMux I__3657 (
            .O(N__18568),
            .I(N__18554));
    Span4Mux_h I__3656 (
            .O(N__18565),
            .I(N__18551));
    InMux I__3655 (
            .O(N__18564),
            .I(N__18546));
    InMux I__3654 (
            .O(N__18563),
            .I(N__18546));
    Span4Mux_h I__3653 (
            .O(N__18560),
            .I(N__18541));
    LocalMux I__3652 (
            .O(N__18557),
            .I(N__18541));
    LocalMux I__3651 (
            .O(N__18554),
            .I(\spi_slave_1.bitcnt_txZ0Z_4 ));
    Odrv4 I__3650 (
            .O(N__18551),
            .I(\spi_slave_1.bitcnt_txZ0Z_4 ));
    LocalMux I__3649 (
            .O(N__18546),
            .I(\spi_slave_1.bitcnt_txZ0Z_4 ));
    Odrv4 I__3648 (
            .O(N__18541),
            .I(\spi_slave_1.bitcnt_txZ0Z_4 ));
    InMux I__3647 (
            .O(N__18532),
            .I(N__18523));
    InMux I__3646 (
            .O(N__18531),
            .I(N__18523));
    InMux I__3645 (
            .O(N__18530),
            .I(N__18523));
    LocalMux I__3644 (
            .O(N__18523),
            .I(N__18518));
    InMux I__3643 (
            .O(N__18522),
            .I(N__18513));
    InMux I__3642 (
            .O(N__18521),
            .I(N__18513));
    Span4Mux_h I__3641 (
            .O(N__18518),
            .I(N__18499));
    LocalMux I__3640 (
            .O(N__18513),
            .I(N__18499));
    InMux I__3639 (
            .O(N__18512),
            .I(N__18496));
    InMux I__3638 (
            .O(N__18511),
            .I(N__18493));
    InMux I__3637 (
            .O(N__18510),
            .I(N__18486));
    InMux I__3636 (
            .O(N__18509),
            .I(N__18486));
    InMux I__3635 (
            .O(N__18508),
            .I(N__18486));
    InMux I__3634 (
            .O(N__18507),
            .I(N__18477));
    InMux I__3633 (
            .O(N__18506),
            .I(N__18477));
    InMux I__3632 (
            .O(N__18505),
            .I(N__18477));
    InMux I__3631 (
            .O(N__18504),
            .I(N__18477));
    Span4Mux_h I__3630 (
            .O(N__18499),
            .I(N__18474));
    LocalMux I__3629 (
            .O(N__18496),
            .I(\spi_slave_1.bitcnt_txZ0Z_0 ));
    LocalMux I__3628 (
            .O(N__18493),
            .I(\spi_slave_1.bitcnt_txZ0Z_0 ));
    LocalMux I__3627 (
            .O(N__18486),
            .I(\spi_slave_1.bitcnt_txZ0Z_0 ));
    LocalMux I__3626 (
            .O(N__18477),
            .I(\spi_slave_1.bitcnt_txZ0Z_0 ));
    Odrv4 I__3625 (
            .O(N__18474),
            .I(\spi_slave_1.bitcnt_txZ0Z_0 ));
    CascadeMux I__3624 (
            .O(N__18463),
            .I(\spi_slave_1.N_58_0_cascade_ ));
    InMux I__3623 (
            .O(N__18460),
            .I(N__18457));
    LocalMux I__3622 (
            .O(N__18457),
            .I(\spi_slave_1.miso_data_outZ0Z_15 ));
    InMux I__3621 (
            .O(N__18454),
            .I(N__18451));
    LocalMux I__3620 (
            .O(N__18451),
            .I(N__18448));
    Span4Mux_h I__3619 (
            .O(N__18448),
            .I(N__18445));
    Odrv4 I__3618 (
            .O(N__18445),
            .I(\spi_slave_1.N_55_0 ));
    InMux I__3617 (
            .O(N__18442),
            .I(N__18439));
    LocalMux I__3616 (
            .O(N__18439),
            .I(N__18435));
    InMux I__3615 (
            .O(N__18438),
            .I(N__18432));
    Odrv4 I__3614 (
            .O(N__18435),
            .I(\spi_slave_1.mosi_data_inZ0Z_15 ));
    LocalMux I__3613 (
            .O(N__18432),
            .I(\spi_slave_1.mosi_data_inZ0Z_15 ));
    CEMux I__3612 (
            .O(N__18427),
            .I(N__18415));
    CEMux I__3611 (
            .O(N__18426),
            .I(N__18415));
    CEMux I__3610 (
            .O(N__18425),
            .I(N__18415));
    CEMux I__3609 (
            .O(N__18424),
            .I(N__18415));
    GlobalMux I__3608 (
            .O(N__18415),
            .I(N__18412));
    gio2CtrlBuf I__3607 (
            .O(N__18412),
            .I(\spi_slave_1.un3_mosi_data_out_g ));
    CascadeMux I__3606 (
            .O(N__18409),
            .I(\sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_ ));
    InMux I__3605 (
            .O(N__18406),
            .I(N__18393));
    InMux I__3604 (
            .O(N__18405),
            .I(N__18393));
    InMux I__3603 (
            .O(N__18404),
            .I(N__18393));
    InMux I__3602 (
            .O(N__18403),
            .I(N__18393));
    CascadeMux I__3601 (
            .O(N__18402),
            .I(N__18389));
    LocalMux I__3600 (
            .O(N__18393),
            .I(N__18386));
    InMux I__3599 (
            .O(N__18392),
            .I(N__18381));
    InMux I__3598 (
            .O(N__18389),
            .I(N__18381));
    Odrv4 I__3597 (
            .O(N__18386),
            .I(\sb_translator_1.num_ledsZ0Z_5 ));
    LocalMux I__3596 (
            .O(N__18381),
            .I(\sb_translator_1.num_ledsZ0Z_5 ));
    CascadeMux I__3595 (
            .O(N__18376),
            .I(\sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_ ));
    InMux I__3594 (
            .O(N__18373),
            .I(N__18368));
    InMux I__3593 (
            .O(N__18372),
            .I(N__18363));
    InMux I__3592 (
            .O(N__18371),
            .I(N__18363));
    LocalMux I__3591 (
            .O(N__18368),
            .I(\demux.N_239 ));
    LocalMux I__3590 (
            .O(N__18363),
            .I(\demux.N_239 ));
    InMux I__3589 (
            .O(N__18358),
            .I(N__18353));
    InMux I__3588 (
            .O(N__18357),
            .I(N__18348));
    InMux I__3587 (
            .O(N__18356),
            .I(N__18348));
    LocalMux I__3586 (
            .O(N__18353),
            .I(\demux.N_241 ));
    LocalMux I__3585 (
            .O(N__18348),
            .I(\demux.N_241 ));
    InMux I__3584 (
            .O(N__18343),
            .I(N__18336));
    InMux I__3583 (
            .O(N__18342),
            .I(N__18336));
    InMux I__3582 (
            .O(N__18341),
            .I(N__18333));
    LocalMux I__3581 (
            .O(N__18336),
            .I(\demux.N_915 ));
    LocalMux I__3580 (
            .O(N__18333),
            .I(\demux.N_915 ));
    CascadeMux I__3579 (
            .O(N__18328),
            .I(N__18325));
    InMux I__3578 (
            .O(N__18325),
            .I(N__18317));
    InMux I__3577 (
            .O(N__18324),
            .I(N__18317));
    InMux I__3576 (
            .O(N__18323),
            .I(N__18312));
    InMux I__3575 (
            .O(N__18322),
            .I(N__18312));
    LocalMux I__3574 (
            .O(N__18317),
            .I(ram_sel_12));
    LocalMux I__3573 (
            .O(N__18312),
            .I(ram_sel_12));
    CascadeMux I__3572 (
            .O(N__18307),
            .I(\demux.N_915_cascade_ ));
    InMux I__3571 (
            .O(N__18304),
            .I(N__18296));
    InMux I__3570 (
            .O(N__18303),
            .I(N__18296));
    InMux I__3569 (
            .O(N__18302),
            .I(N__18291));
    InMux I__3568 (
            .O(N__18301),
            .I(N__18291));
    LocalMux I__3567 (
            .O(N__18296),
            .I(ram_sel_2));
    LocalMux I__3566 (
            .O(N__18291),
            .I(ram_sel_2));
    InMux I__3565 (
            .O(N__18286),
            .I(N__18281));
    CascadeMux I__3564 (
            .O(N__18285),
            .I(N__18278));
    CascadeMux I__3563 (
            .O(N__18284),
            .I(N__18275));
    LocalMux I__3562 (
            .O(N__18281),
            .I(N__18270));
    InMux I__3561 (
            .O(N__18278),
            .I(N__18263));
    InMux I__3560 (
            .O(N__18275),
            .I(N__18263));
    InMux I__3559 (
            .O(N__18274),
            .I(N__18263));
    InMux I__3558 (
            .O(N__18273),
            .I(N__18260));
    Odrv4 I__3557 (
            .O(N__18270),
            .I(ram_sel_3));
    LocalMux I__3556 (
            .O(N__18263),
            .I(ram_sel_3));
    LocalMux I__3555 (
            .O(N__18260),
            .I(ram_sel_3));
    CascadeMux I__3554 (
            .O(N__18253),
            .I(N__18247));
    InMux I__3553 (
            .O(N__18252),
            .I(N__18239));
    InMux I__3552 (
            .O(N__18251),
            .I(N__18239));
    InMux I__3551 (
            .O(N__18250),
            .I(N__18239));
    InMux I__3550 (
            .O(N__18247),
            .I(N__18234));
    InMux I__3549 (
            .O(N__18246),
            .I(N__18234));
    LocalMux I__3548 (
            .O(N__18239),
            .I(ram_sel_8));
    LocalMux I__3547 (
            .O(N__18234),
            .I(ram_sel_8));
    CascadeMux I__3546 (
            .O(N__18229),
            .I(N__18223));
    CascadeMux I__3545 (
            .O(N__18228),
            .I(N__18220));
    CascadeMux I__3544 (
            .O(N__18227),
            .I(N__18217));
    CascadeMux I__3543 (
            .O(N__18226),
            .I(N__18214));
    CascadeBuf I__3542 (
            .O(N__18223),
            .I(N__18211));
    CascadeBuf I__3541 (
            .O(N__18220),
            .I(N__18208));
    CascadeBuf I__3540 (
            .O(N__18217),
            .I(N__18205));
    CascadeBuf I__3539 (
            .O(N__18214),
            .I(N__18202));
    CascadeMux I__3538 (
            .O(N__18211),
            .I(N__18199));
    CascadeMux I__3537 (
            .O(N__18208),
            .I(N__18196));
    CascadeMux I__3536 (
            .O(N__18205),
            .I(N__18193));
    CascadeMux I__3535 (
            .O(N__18202),
            .I(N__18190));
    CascadeBuf I__3534 (
            .O(N__18199),
            .I(N__18187));
    CascadeBuf I__3533 (
            .O(N__18196),
            .I(N__18184));
    CascadeBuf I__3532 (
            .O(N__18193),
            .I(N__18181));
    CascadeBuf I__3531 (
            .O(N__18190),
            .I(N__18178));
    CascadeMux I__3530 (
            .O(N__18187),
            .I(N__18175));
    CascadeMux I__3529 (
            .O(N__18184),
            .I(N__18172));
    CascadeMux I__3528 (
            .O(N__18181),
            .I(N__18169));
    CascadeMux I__3527 (
            .O(N__18178),
            .I(N__18166));
    CascadeBuf I__3526 (
            .O(N__18175),
            .I(N__18163));
    CascadeBuf I__3525 (
            .O(N__18172),
            .I(N__18160));
    CascadeBuf I__3524 (
            .O(N__18169),
            .I(N__18157));
    CascadeBuf I__3523 (
            .O(N__18166),
            .I(N__18154));
    CascadeMux I__3522 (
            .O(N__18163),
            .I(N__18151));
    CascadeMux I__3521 (
            .O(N__18160),
            .I(N__18148));
    CascadeMux I__3520 (
            .O(N__18157),
            .I(N__18145));
    CascadeMux I__3519 (
            .O(N__18154),
            .I(N__18142));
    CascadeBuf I__3518 (
            .O(N__18151),
            .I(N__18139));
    CascadeBuf I__3517 (
            .O(N__18148),
            .I(N__18136));
    CascadeBuf I__3516 (
            .O(N__18145),
            .I(N__18133));
    CascadeBuf I__3515 (
            .O(N__18142),
            .I(N__18130));
    CascadeMux I__3514 (
            .O(N__18139),
            .I(N__18127));
    CascadeMux I__3513 (
            .O(N__18136),
            .I(N__18124));
    CascadeMux I__3512 (
            .O(N__18133),
            .I(N__18121));
    CascadeMux I__3511 (
            .O(N__18130),
            .I(N__18118));
    CascadeBuf I__3510 (
            .O(N__18127),
            .I(N__18115));
    CascadeBuf I__3509 (
            .O(N__18124),
            .I(N__18112));
    CascadeBuf I__3508 (
            .O(N__18121),
            .I(N__18109));
    CascadeBuf I__3507 (
            .O(N__18118),
            .I(N__18106));
    CascadeMux I__3506 (
            .O(N__18115),
            .I(N__18103));
    CascadeMux I__3505 (
            .O(N__18112),
            .I(N__18100));
    CascadeMux I__3504 (
            .O(N__18109),
            .I(N__18097));
    CascadeMux I__3503 (
            .O(N__18106),
            .I(N__18094));
    CascadeBuf I__3502 (
            .O(N__18103),
            .I(N__18091));
    CascadeBuf I__3501 (
            .O(N__18100),
            .I(N__18088));
    CascadeBuf I__3500 (
            .O(N__18097),
            .I(N__18085));
    CascadeBuf I__3499 (
            .O(N__18094),
            .I(N__18082));
    CascadeMux I__3498 (
            .O(N__18091),
            .I(N__18079));
    CascadeMux I__3497 (
            .O(N__18088),
            .I(N__18076));
    CascadeMux I__3496 (
            .O(N__18085),
            .I(N__18073));
    CascadeMux I__3495 (
            .O(N__18082),
            .I(N__18070));
    InMux I__3494 (
            .O(N__18079),
            .I(N__18067));
    InMux I__3493 (
            .O(N__18076),
            .I(N__18064));
    InMux I__3492 (
            .O(N__18073),
            .I(N__18061));
    InMux I__3491 (
            .O(N__18070),
            .I(N__18058));
    LocalMux I__3490 (
            .O(N__18067),
            .I(N__18052));
    LocalMux I__3489 (
            .O(N__18064),
            .I(N__18052));
    LocalMux I__3488 (
            .O(N__18061),
            .I(N__18047));
    LocalMux I__3487 (
            .O(N__18058),
            .I(N__18047));
    InMux I__3486 (
            .O(N__18057),
            .I(N__18044));
    Span4Mux_s2_v I__3485 (
            .O(N__18052),
            .I(N__18041));
    Span4Mux_s2_v I__3484 (
            .O(N__18047),
            .I(N__18038));
    LocalMux I__3483 (
            .O(N__18044),
            .I(addr_out_8));
    Odrv4 I__3482 (
            .O(N__18041),
            .I(addr_out_8));
    Odrv4 I__3481 (
            .O(N__18038),
            .I(addr_out_8));
    CEMux I__3480 (
            .O(N__18031),
            .I(N__18028));
    LocalMux I__3479 (
            .O(N__18028),
            .I(N__18024));
    CEMux I__3478 (
            .O(N__18027),
            .I(N__18021));
    Span4Mux_v I__3477 (
            .O(N__18024),
            .I(N__18018));
    LocalMux I__3476 (
            .O(N__18021),
            .I(N__18015));
    Odrv4 I__3475 (
            .O(N__18018),
            .I(\sb_translator_1.state_RNI88IGAZ0Z_0 ));
    Odrv12 I__3474 (
            .O(N__18015),
            .I(\sb_translator_1.state_RNI88IGAZ0Z_0 ));
    IoInMux I__3473 (
            .O(N__18010),
            .I(N__18007));
    LocalMux I__3472 (
            .O(N__18007),
            .I(N__18004));
    Span4Mux_s0_v I__3471 (
            .O(N__18004),
            .I(N__18001));
    Odrv4 I__3470 (
            .O(N__18001),
            .I(\sb_translator_1.state_leds_2_sqmuxa ));
    CascadeMux I__3469 (
            .O(N__17998),
            .I(N__17994));
    CascadeMux I__3468 (
            .O(N__17997),
            .I(N__17990));
    InMux I__3467 (
            .O(N__17994),
            .I(N__17985));
    InMux I__3466 (
            .O(N__17993),
            .I(N__17985));
    InMux I__3465 (
            .O(N__17990),
            .I(N__17982));
    LocalMux I__3464 (
            .O(N__17985),
            .I(N__17979));
    LocalMux I__3463 (
            .O(N__17982),
            .I(\sb_translator_1.state_ledsZ0 ));
    Odrv12 I__3462 (
            .O(N__17979),
            .I(\sb_translator_1.state_ledsZ0 ));
    InMux I__3461 (
            .O(N__17974),
            .I(N__17971));
    LocalMux I__3460 (
            .O(N__17971),
            .I(\spi_slave_1.miso_data_outZ0Z_9 ));
    InMux I__3459 (
            .O(N__17968),
            .I(N__17965));
    LocalMux I__3458 (
            .O(N__17965),
            .I(\spi_slave_1.miso_data_outZ0Z_10 ));
    InMux I__3457 (
            .O(N__17962),
            .I(N__17959));
    LocalMux I__3456 (
            .O(N__17959),
            .I(N__17956));
    Odrv4 I__3455 (
            .O(N__17956),
            .I(\spi_slave_1.miso_RNOZ0Z_13 ));
    CascadeMux I__3454 (
            .O(N__17953),
            .I(\demux.N_242_cascade_ ));
    CascadeMux I__3453 (
            .O(N__17950),
            .I(\demux.N_424_i_0_a2Z0Z_34_cascade_ ));
    InMux I__3452 (
            .O(N__17947),
            .I(N__17938));
    InMux I__3451 (
            .O(N__17946),
            .I(N__17938));
    InMux I__3450 (
            .O(N__17945),
            .I(N__17928));
    InMux I__3449 (
            .O(N__17944),
            .I(N__17928));
    InMux I__3448 (
            .O(N__17943),
            .I(N__17928));
    LocalMux I__3447 (
            .O(N__17938),
            .I(N__17925));
    InMux I__3446 (
            .O(N__17937),
            .I(N__17918));
    InMux I__3445 (
            .O(N__17936),
            .I(N__17918));
    InMux I__3444 (
            .O(N__17935),
            .I(N__17918));
    LocalMux I__3443 (
            .O(N__17928),
            .I(N__17915));
    Span4Mux_h I__3442 (
            .O(N__17925),
            .I(N__17912));
    LocalMux I__3441 (
            .O(N__17918),
            .I(\demux.N_424_i_0_aZ0Z2 ));
    Odrv4 I__3440 (
            .O(N__17915),
            .I(\demux.N_424_i_0_aZ0Z2 ));
    Odrv4 I__3439 (
            .O(N__17912),
            .I(\demux.N_424_i_0_aZ0Z2 ));
    InMux I__3438 (
            .O(N__17905),
            .I(N__17901));
    InMux I__3437 (
            .O(N__17904),
            .I(N__17898));
    LocalMux I__3436 (
            .O(N__17901),
            .I(\demux.N_242 ));
    LocalMux I__3435 (
            .O(N__17898),
            .I(\demux.N_242 ));
    InMux I__3434 (
            .O(N__17893),
            .I(N__17884));
    InMux I__3433 (
            .O(N__17892),
            .I(N__17884));
    InMux I__3432 (
            .O(N__17891),
            .I(N__17884));
    LocalMux I__3431 (
            .O(N__17884),
            .I(\demux.N_916 ));
    CascadeMux I__3430 (
            .O(N__17881),
            .I(N__17876));
    InMux I__3429 (
            .O(N__17880),
            .I(N__17872));
    InMux I__3428 (
            .O(N__17879),
            .I(N__17865));
    InMux I__3427 (
            .O(N__17876),
            .I(N__17865));
    InMux I__3426 (
            .O(N__17875),
            .I(N__17865));
    LocalMux I__3425 (
            .O(N__17872),
            .I(ram_sel_5));
    LocalMux I__3424 (
            .O(N__17865),
            .I(ram_sel_5));
    CascadeMux I__3423 (
            .O(N__17860),
            .I(\demux.N_916_cascade_ ));
    InMux I__3422 (
            .O(N__17857),
            .I(N__17851));
    InMux I__3421 (
            .O(N__17856),
            .I(N__17848));
    InMux I__3420 (
            .O(N__17855),
            .I(N__17843));
    InMux I__3419 (
            .O(N__17854),
            .I(N__17843));
    LocalMux I__3418 (
            .O(N__17851),
            .I(ram_sel_1));
    LocalMux I__3417 (
            .O(N__17848),
            .I(ram_sel_1));
    LocalMux I__3416 (
            .O(N__17843),
            .I(ram_sel_1));
    CascadeMux I__3415 (
            .O(N__17836),
            .I(\sb_translator_1.num_leds_1_sqmuxa_cascade_ ));
    InMux I__3414 (
            .O(N__17833),
            .I(N__17826));
    InMux I__3413 (
            .O(N__17832),
            .I(N__17826));
    InMux I__3412 (
            .O(N__17831),
            .I(N__17823));
    LocalMux I__3411 (
            .O(N__17826),
            .I(N__17818));
    LocalMux I__3410 (
            .O(N__17823),
            .I(N__17818));
    Span4Mux_v I__3409 (
            .O(N__17818),
            .I(N__17815));
    Odrv4 I__3408 (
            .O(N__17815),
            .I(\sb_translator_1.send_leds_n_1_sqmuxa ));
    InMux I__3407 (
            .O(N__17812),
            .I(N__17809));
    LocalMux I__3406 (
            .O(N__17809),
            .I(\sb_translator_1.N_59 ));
    InMux I__3405 (
            .O(N__17806),
            .I(N__17803));
    LocalMux I__3404 (
            .O(N__17803),
            .I(N__17800));
    Span4Mux_h I__3403 (
            .O(N__17800),
            .I(N__17797));
    Odrv4 I__3402 (
            .O(N__17797),
            .I(miso_data_in_0));
    InMux I__3401 (
            .O(N__17794),
            .I(N__17789));
    CascadeMux I__3400 (
            .O(N__17793),
            .I(N__17785));
    InMux I__3399 (
            .O(N__17792),
            .I(N__17782));
    LocalMux I__3398 (
            .O(N__17789),
            .I(N__17779));
    InMux I__3397 (
            .O(N__17788),
            .I(N__17774));
    InMux I__3396 (
            .O(N__17785),
            .I(N__17774));
    LocalMux I__3395 (
            .O(N__17782),
            .I(N__17771));
    Span4Mux_v I__3394 (
            .O(N__17779),
            .I(N__17768));
    LocalMux I__3393 (
            .O(N__17774),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5 ));
    Odrv4 I__3392 (
            .O(N__17771),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5 ));
    Odrv4 I__3391 (
            .O(N__17768),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5 ));
    InMux I__3390 (
            .O(N__17761),
            .I(N__17758));
    LocalMux I__3389 (
            .O(N__17758),
            .I(N__17754));
    InMux I__3388 (
            .O(N__17757),
            .I(N__17751));
    Span4Mux_v I__3387 (
            .O(N__17754),
            .I(N__17746));
    LocalMux I__3386 (
            .O(N__17751),
            .I(N__17743));
    InMux I__3385 (
            .O(N__17750),
            .I(N__17740));
    InMux I__3384 (
            .O(N__17749),
            .I(N__17737));
    Odrv4 I__3383 (
            .O(N__17746),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ));
    Odrv4 I__3382 (
            .O(N__17743),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ));
    LocalMux I__3381 (
            .O(N__17740),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ));
    LocalMux I__3380 (
            .O(N__17737),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ));
    CascadeMux I__3379 (
            .O(N__17728),
            .I(N__17724));
    InMux I__3378 (
            .O(N__17727),
            .I(N__17721));
    InMux I__3377 (
            .O(N__17724),
            .I(N__17716));
    LocalMux I__3376 (
            .O(N__17721),
            .I(N__17713));
    InMux I__3375 (
            .O(N__17720),
            .I(N__17708));
    InMux I__3374 (
            .O(N__17719),
            .I(N__17708));
    LocalMux I__3373 (
            .O(N__17716),
            .I(N__17705));
    Span4Mux_v I__3372 (
            .O(N__17713),
            .I(N__17702));
    LocalMux I__3371 (
            .O(N__17708),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0 ));
    Odrv4 I__3370 (
            .O(N__17705),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0 ));
    Odrv4 I__3369 (
            .O(N__17702),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0 ));
    InMux I__3368 (
            .O(N__17695),
            .I(N__17683));
    InMux I__3367 (
            .O(N__17694),
            .I(N__17683));
    InMux I__3366 (
            .O(N__17693),
            .I(N__17683));
    InMux I__3365 (
            .O(N__17692),
            .I(N__17683));
    LocalMux I__3364 (
            .O(N__17683),
            .I(N__17676));
    InMux I__3363 (
            .O(N__17682),
            .I(N__17671));
    InMux I__3362 (
            .O(N__17681),
            .I(N__17671));
    InMux I__3361 (
            .O(N__17680),
            .I(N__17668));
    InMux I__3360 (
            .O(N__17679),
            .I(N__17665));
    Span4Mux_v I__3359 (
            .O(N__17676),
            .I(N__17660));
    LocalMux I__3358 (
            .O(N__17671),
            .I(N__17660));
    LocalMux I__3357 (
            .O(N__17668),
            .I(N__17655));
    LocalMux I__3356 (
            .O(N__17665),
            .I(N__17655));
    Span4Mux_v I__3355 (
            .O(N__17660),
            .I(N__17652));
    Span4Mux_v I__3354 (
            .O(N__17655),
            .I(N__17649));
    Odrv4 I__3353 (
            .O(N__17652),
            .I(mosi_data_out_18));
    Odrv4 I__3352 (
            .O(N__17649),
            .I(mosi_data_out_18));
    InMux I__3351 (
            .O(N__17644),
            .I(N__17636));
    InMux I__3350 (
            .O(N__17643),
            .I(N__17636));
    InMux I__3349 (
            .O(N__17642),
            .I(N__17631));
    InMux I__3348 (
            .O(N__17641),
            .I(N__17631));
    LocalMux I__3347 (
            .O(N__17636),
            .I(N__17624));
    LocalMux I__3346 (
            .O(N__17631),
            .I(N__17624));
    InMux I__3345 (
            .O(N__17630),
            .I(N__17617));
    InMux I__3344 (
            .O(N__17629),
            .I(N__17617));
    Span4Mux_v I__3343 (
            .O(N__17624),
            .I(N__17614));
    InMux I__3342 (
            .O(N__17623),
            .I(N__17609));
    InMux I__3341 (
            .O(N__17622),
            .I(N__17609));
    LocalMux I__3340 (
            .O(N__17617),
            .I(N__17606));
    Span4Mux_h I__3339 (
            .O(N__17614),
            .I(N__17601));
    LocalMux I__3338 (
            .O(N__17609),
            .I(N__17601));
    Span12Mux_s11_h I__3337 (
            .O(N__17606),
            .I(N__17598));
    Span4Mux_v I__3336 (
            .O(N__17601),
            .I(N__17595));
    Odrv12 I__3335 (
            .O(N__17598),
            .I(mosi_data_out_19));
    Odrv4 I__3334 (
            .O(N__17595),
            .I(mosi_data_out_19));
    InMux I__3333 (
            .O(N__17590),
            .I(N__17578));
    InMux I__3332 (
            .O(N__17589),
            .I(N__17578));
    InMux I__3331 (
            .O(N__17588),
            .I(N__17578));
    InMux I__3330 (
            .O(N__17587),
            .I(N__17578));
    LocalMux I__3329 (
            .O(N__17578),
            .I(N__17573));
    InMux I__3328 (
            .O(N__17577),
            .I(N__17568));
    InMux I__3327 (
            .O(N__17576),
            .I(N__17565));
    Span4Mux_v I__3326 (
            .O(N__17573),
            .I(N__17562));
    InMux I__3325 (
            .O(N__17572),
            .I(N__17557));
    InMux I__3324 (
            .O(N__17571),
            .I(N__17557));
    LocalMux I__3323 (
            .O(N__17568),
            .I(N__17552));
    LocalMux I__3322 (
            .O(N__17565),
            .I(N__17552));
    Span4Mux_h I__3321 (
            .O(N__17562),
            .I(N__17547));
    LocalMux I__3320 (
            .O(N__17557),
            .I(N__17547));
    Span4Mux_v I__3319 (
            .O(N__17552),
            .I(N__17544));
    Span4Mux_v I__3318 (
            .O(N__17547),
            .I(N__17541));
    Odrv4 I__3317 (
            .O(N__17544),
            .I(mosi_data_out_20));
    Odrv4 I__3316 (
            .O(N__17541),
            .I(mosi_data_out_20));
    CascadeMux I__3315 (
            .O(N__17536),
            .I(N__17533));
    InMux I__3314 (
            .O(N__17533),
            .I(N__17530));
    LocalMux I__3313 (
            .O(N__17530),
            .I(N__17524));
    InMux I__3312 (
            .O(N__17529),
            .I(N__17521));
    CascadeMux I__3311 (
            .O(N__17528),
            .I(N__17518));
    CascadeMux I__3310 (
            .O(N__17527),
            .I(N__17515));
    Span4Mux_v I__3309 (
            .O(N__17524),
            .I(N__17512));
    LocalMux I__3308 (
            .O(N__17521),
            .I(N__17509));
    InMux I__3307 (
            .O(N__17518),
            .I(N__17504));
    InMux I__3306 (
            .O(N__17515),
            .I(N__17504));
    Odrv4 I__3305 (
            .O(N__17512),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3 ));
    Odrv4 I__3304 (
            .O(N__17509),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3 ));
    LocalMux I__3303 (
            .O(N__17504),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3 ));
    CascadeMux I__3302 (
            .O(N__17497),
            .I(\demux.N_238_cascade_ ));
    CEMux I__3301 (
            .O(N__17494),
            .I(N__17490));
    InMux I__3300 (
            .O(N__17493),
            .I(N__17487));
    LocalMux I__3299 (
            .O(N__17490),
            .I(N__17484));
    LocalMux I__3298 (
            .O(N__17487),
            .I(N__17479));
    Span4Mux_v I__3297 (
            .O(N__17484),
            .I(N__17476));
    CEMux I__3296 (
            .O(N__17483),
            .I(N__17473));
    CEMux I__3295 (
            .O(N__17482),
            .I(N__17470));
    Span12Mux_s9_h I__3294 (
            .O(N__17479),
            .I(N__17467));
    Odrv4 I__3293 (
            .O(N__17476),
            .I(\sb_translator_1.N_58 ));
    LocalMux I__3292 (
            .O(N__17473),
            .I(\sb_translator_1.N_58 ));
    LocalMux I__3291 (
            .O(N__17470),
            .I(\sb_translator_1.N_58 ));
    Odrv12 I__3290 (
            .O(N__17467),
            .I(\sb_translator_1.N_58 ));
    InMux I__3289 (
            .O(N__17458),
            .I(N__17455));
    LocalMux I__3288 (
            .O(N__17455),
            .I(\sb_translator_1.state_RNIEL0N9_0Z0Z_6 ));
    CascadeMux I__3287 (
            .O(N__17452),
            .I(N__17444));
    InMux I__3286 (
            .O(N__17451),
            .I(N__17432));
    InMux I__3285 (
            .O(N__17450),
            .I(N__17432));
    InMux I__3284 (
            .O(N__17449),
            .I(N__17432));
    InMux I__3283 (
            .O(N__17448),
            .I(N__17432));
    InMux I__3282 (
            .O(N__17447),
            .I(N__17432));
    InMux I__3281 (
            .O(N__17444),
            .I(N__17427));
    InMux I__3280 (
            .O(N__17443),
            .I(N__17427));
    LocalMux I__3279 (
            .O(N__17432),
            .I(N__17424));
    LocalMux I__3278 (
            .O(N__17427),
            .I(\sb_translator_1.cnt_ram_readZ0Z_0 ));
    Odrv12 I__3277 (
            .O(N__17424),
            .I(\sb_translator_1.cnt_ram_readZ0Z_0 ));
    CascadeMux I__3276 (
            .O(N__17419),
            .I(N__17413));
    CascadeMux I__3275 (
            .O(N__17418),
            .I(N__17410));
    CascadeMux I__3274 (
            .O(N__17417),
            .I(N__17407));
    CascadeMux I__3273 (
            .O(N__17416),
            .I(N__17403));
    InMux I__3272 (
            .O(N__17413),
            .I(N__17399));
    InMux I__3271 (
            .O(N__17410),
            .I(N__17388));
    InMux I__3270 (
            .O(N__17407),
            .I(N__17388));
    InMux I__3269 (
            .O(N__17406),
            .I(N__17388));
    InMux I__3268 (
            .O(N__17403),
            .I(N__17388));
    InMux I__3267 (
            .O(N__17402),
            .I(N__17388));
    LocalMux I__3266 (
            .O(N__17399),
            .I(N__17383));
    LocalMux I__3265 (
            .O(N__17388),
            .I(N__17383));
    Odrv12 I__3264 (
            .O(N__17383),
            .I(\sb_translator_1.cnt_ram_readZ0Z_1 ));
    InMux I__3263 (
            .O(N__17380),
            .I(N__17377));
    LocalMux I__3262 (
            .O(N__17377),
            .I(N__17374));
    Span4Mux_v I__3261 (
            .O(N__17374),
            .I(N__17371));
    Odrv4 I__3260 (
            .O(N__17371),
            .I(demux_data_in_42));
    InMux I__3259 (
            .O(N__17368),
            .I(N__17364));
    InMux I__3258 (
            .O(N__17367),
            .I(N__17361));
    LocalMux I__3257 (
            .O(N__17364),
            .I(N__17355));
    LocalMux I__3256 (
            .O(N__17361),
            .I(N__17352));
    InMux I__3255 (
            .O(N__17360),
            .I(N__17347));
    InMux I__3254 (
            .O(N__17359),
            .I(N__17347));
    InMux I__3253 (
            .O(N__17358),
            .I(N__17343));
    Span4Mux_v I__3252 (
            .O(N__17355),
            .I(N__17338));
    Span4Mux_v I__3251 (
            .O(N__17352),
            .I(N__17338));
    LocalMux I__3250 (
            .O(N__17347),
            .I(N__17335));
    InMux I__3249 (
            .O(N__17346),
            .I(N__17332));
    LocalMux I__3248 (
            .O(N__17343),
            .I(N__17329));
    Odrv4 I__3247 (
            .O(N__17338),
            .I(\sb_translator_1.cntZ0Z_11 ));
    Odrv4 I__3246 (
            .O(N__17335),
            .I(\sb_translator_1.cntZ0Z_11 ));
    LocalMux I__3245 (
            .O(N__17332),
            .I(\sb_translator_1.cntZ0Z_11 ));
    Odrv4 I__3244 (
            .O(N__17329),
            .I(\sb_translator_1.cntZ0Z_11 ));
    InMux I__3243 (
            .O(N__17320),
            .I(N__17316));
    InMux I__3242 (
            .O(N__17319),
            .I(N__17313));
    LocalMux I__3241 (
            .O(N__17316),
            .I(N__17308));
    LocalMux I__3240 (
            .O(N__17313),
            .I(N__17305));
    InMux I__3239 (
            .O(N__17312),
            .I(N__17300));
    InMux I__3238 (
            .O(N__17311),
            .I(N__17300));
    Span4Mux_v I__3237 (
            .O(N__17308),
            .I(N__17293));
    Span4Mux_v I__3236 (
            .O(N__17305),
            .I(N__17293));
    LocalMux I__3235 (
            .O(N__17300),
            .I(N__17293));
    Span4Mux_h I__3234 (
            .O(N__17293),
            .I(N__17288));
    InMux I__3233 (
            .O(N__17292),
            .I(N__17285));
    InMux I__3232 (
            .O(N__17291),
            .I(N__17282));
    Odrv4 I__3231 (
            .O(N__17288),
            .I(\sb_translator_1.cntZ0Z_10 ));
    LocalMux I__3230 (
            .O(N__17285),
            .I(\sb_translator_1.cntZ0Z_10 ));
    LocalMux I__3229 (
            .O(N__17282),
            .I(\sb_translator_1.cntZ0Z_10 ));
    CascadeMux I__3228 (
            .O(N__17275),
            .I(N__17272));
    InMux I__3227 (
            .O(N__17272),
            .I(N__17269));
    LocalMux I__3226 (
            .O(N__17269),
            .I(N__17266));
    Span4Mux_v I__3225 (
            .O(N__17266),
            .I(N__17262));
    CascadeMux I__3224 (
            .O(N__17265),
            .I(N__17259));
    Span4Mux_h I__3223 (
            .O(N__17262),
            .I(N__17256));
    InMux I__3222 (
            .O(N__17259),
            .I(N__17253));
    Odrv4 I__3221 (
            .O(N__17256),
            .I(\sb_translator_1.ram_we_6_0_0_a2_0_6 ));
    LocalMux I__3220 (
            .O(N__17253),
            .I(\sb_translator_1.ram_we_6_0_0_a2_0_6 ));
    InMux I__3219 (
            .O(N__17248),
            .I(N__17245));
    LocalMux I__3218 (
            .O(N__17245),
            .I(N__17242));
    Span4Mux_v I__3217 (
            .O(N__17242),
            .I(N__17239));
    Odrv4 I__3216 (
            .O(N__17239),
            .I(miso_data_in_2));
    CascadeMux I__3215 (
            .O(N__17236),
            .I(N__17229));
    InMux I__3214 (
            .O(N__17235),
            .I(N__17224));
    CascadeMux I__3213 (
            .O(N__17234),
            .I(N__17217));
    InMux I__3212 (
            .O(N__17233),
            .I(N__17210));
    InMux I__3211 (
            .O(N__17232),
            .I(N__17210));
    InMux I__3210 (
            .O(N__17229),
            .I(N__17210));
    CascadeMux I__3209 (
            .O(N__17228),
            .I(N__17207));
    CascadeMux I__3208 (
            .O(N__17227),
            .I(N__17204));
    LocalMux I__3207 (
            .O(N__17224),
            .I(N__17193));
    CascadeMux I__3206 (
            .O(N__17223),
            .I(N__17190));
    CascadeMux I__3205 (
            .O(N__17222),
            .I(N__17187));
    CascadeMux I__3204 (
            .O(N__17221),
            .I(N__17184));
    CascadeMux I__3203 (
            .O(N__17220),
            .I(N__17181));
    InMux I__3202 (
            .O(N__17217),
            .I(N__17174));
    LocalMux I__3201 (
            .O(N__17210),
            .I(N__17171));
    InMux I__3200 (
            .O(N__17207),
            .I(N__17164));
    InMux I__3199 (
            .O(N__17204),
            .I(N__17164));
    InMux I__3198 (
            .O(N__17203),
            .I(N__17164));
    InMux I__3197 (
            .O(N__17202),
            .I(N__17149));
    InMux I__3196 (
            .O(N__17201),
            .I(N__17149));
    InMux I__3195 (
            .O(N__17200),
            .I(N__17149));
    InMux I__3194 (
            .O(N__17199),
            .I(N__17149));
    InMux I__3193 (
            .O(N__17198),
            .I(N__17149));
    InMux I__3192 (
            .O(N__17197),
            .I(N__17149));
    InMux I__3191 (
            .O(N__17196),
            .I(N__17149));
    Span4Mux_v I__3190 (
            .O(N__17193),
            .I(N__17146));
    InMux I__3189 (
            .O(N__17190),
            .I(N__17129));
    InMux I__3188 (
            .O(N__17187),
            .I(N__17129));
    InMux I__3187 (
            .O(N__17184),
            .I(N__17129));
    InMux I__3186 (
            .O(N__17181),
            .I(N__17129));
    InMux I__3185 (
            .O(N__17180),
            .I(N__17129));
    InMux I__3184 (
            .O(N__17179),
            .I(N__17129));
    InMux I__3183 (
            .O(N__17178),
            .I(N__17129));
    InMux I__3182 (
            .O(N__17177),
            .I(N__17129));
    LocalMux I__3181 (
            .O(N__17174),
            .I(N__17126));
    Span4Mux_v I__3180 (
            .O(N__17171),
            .I(N__17123));
    LocalMux I__3179 (
            .O(N__17164),
            .I(N__17116));
    LocalMux I__3178 (
            .O(N__17149),
            .I(N__17116));
    Span4Mux_h I__3177 (
            .O(N__17146),
            .I(N__17116));
    LocalMux I__3176 (
            .O(N__17129),
            .I(mosi_data_out_22));
    Odrv4 I__3175 (
            .O(N__17126),
            .I(mosi_data_out_22));
    Odrv4 I__3174 (
            .O(N__17123),
            .I(mosi_data_out_22));
    Odrv4 I__3173 (
            .O(N__17116),
            .I(mosi_data_out_22));
    InMux I__3172 (
            .O(N__17107),
            .I(N__17083));
    InMux I__3171 (
            .O(N__17106),
            .I(N__17083));
    InMux I__3170 (
            .O(N__17105),
            .I(N__17083));
    InMux I__3169 (
            .O(N__17104),
            .I(N__17068));
    InMux I__3168 (
            .O(N__17103),
            .I(N__17068));
    InMux I__3167 (
            .O(N__17102),
            .I(N__17068));
    InMux I__3166 (
            .O(N__17101),
            .I(N__17068));
    InMux I__3165 (
            .O(N__17100),
            .I(N__17068));
    InMux I__3164 (
            .O(N__17099),
            .I(N__17068));
    InMux I__3163 (
            .O(N__17098),
            .I(N__17068));
    InMux I__3162 (
            .O(N__17097),
            .I(N__17051));
    InMux I__3161 (
            .O(N__17096),
            .I(N__17051));
    InMux I__3160 (
            .O(N__17095),
            .I(N__17051));
    InMux I__3159 (
            .O(N__17094),
            .I(N__17051));
    InMux I__3158 (
            .O(N__17093),
            .I(N__17051));
    InMux I__3157 (
            .O(N__17092),
            .I(N__17051));
    InMux I__3156 (
            .O(N__17091),
            .I(N__17051));
    InMux I__3155 (
            .O(N__17090),
            .I(N__17051));
    LocalMux I__3154 (
            .O(N__17083),
            .I(N__17043));
    LocalMux I__3153 (
            .O(N__17068),
            .I(N__17043));
    LocalMux I__3152 (
            .O(N__17051),
            .I(N__17043));
    InMux I__3151 (
            .O(N__17050),
            .I(N__17040));
    Span4Mux_v I__3150 (
            .O(N__17043),
            .I(N__17037));
    LocalMux I__3149 (
            .O(N__17040),
            .I(N__17034));
    Odrv4 I__3148 (
            .O(N__17037),
            .I(\sb_translator_1.N_1087 ));
    Odrv12 I__3147 (
            .O(N__17034),
            .I(\sb_translator_1.N_1087 ));
    InMux I__3146 (
            .O(N__17029),
            .I(N__17026));
    LocalMux I__3145 (
            .O(N__17026),
            .I(N__17021));
    InMux I__3144 (
            .O(N__17025),
            .I(N__17018));
    InMux I__3143 (
            .O(N__17024),
            .I(N__17015));
    Odrv4 I__3142 (
            .O(N__17021),
            .I(mosi_data_out_3));
    LocalMux I__3141 (
            .O(N__17018),
            .I(mosi_data_out_3));
    LocalMux I__3140 (
            .O(N__17015),
            .I(mosi_data_out_3));
    InMux I__3139 (
            .O(N__17008),
            .I(N__17005));
    LocalMux I__3138 (
            .O(N__17005),
            .I(\sb_translator_1.instr_tmpZ1Z_3 ));
    InMux I__3137 (
            .O(N__17002),
            .I(N__16997));
    InMux I__3136 (
            .O(N__17001),
            .I(N__16994));
    InMux I__3135 (
            .O(N__17000),
            .I(N__16991));
    LocalMux I__3134 (
            .O(N__16997),
            .I(N__16988));
    LocalMux I__3133 (
            .O(N__16994),
            .I(mosi_data_out_4));
    LocalMux I__3132 (
            .O(N__16991),
            .I(mosi_data_out_4));
    Odrv12 I__3131 (
            .O(N__16988),
            .I(mosi_data_out_4));
    InMux I__3130 (
            .O(N__16981),
            .I(N__16978));
    LocalMux I__3129 (
            .O(N__16978),
            .I(\sb_translator_1.instr_tmpZ1Z_4 ));
    CEMux I__3128 (
            .O(N__16975),
            .I(N__16972));
    LocalMux I__3127 (
            .O(N__16972),
            .I(N__16968));
    CEMux I__3126 (
            .O(N__16971),
            .I(N__16965));
    Span4Mux_h I__3125 (
            .O(N__16968),
            .I(N__16960));
    LocalMux I__3124 (
            .O(N__16965),
            .I(N__16960));
    Span4Mux_h I__3123 (
            .O(N__16960),
            .I(N__16957));
    Span4Mux_s1_h I__3122 (
            .O(N__16957),
            .I(N__16954));
    Odrv4 I__3121 (
            .O(N__16954),
            .I(\sb_translator_1.state_RNIKJOCZ0Z_5 ));
    InMux I__3120 (
            .O(N__16951),
            .I(N__16947));
    InMux I__3119 (
            .O(N__16950),
            .I(N__16942));
    LocalMux I__3118 (
            .O(N__16947),
            .I(N__16939));
    InMux I__3117 (
            .O(N__16946),
            .I(N__16936));
    InMux I__3116 (
            .O(N__16945),
            .I(N__16933));
    LocalMux I__3115 (
            .O(N__16942),
            .I(N__16930));
    Span4Mux_h I__3114 (
            .O(N__16939),
            .I(N__16927));
    LocalMux I__3113 (
            .O(N__16936),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ));
    LocalMux I__3112 (
            .O(N__16933),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ));
    Odrv12 I__3111 (
            .O(N__16930),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ));
    Odrv4 I__3110 (
            .O(N__16927),
            .I(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ));
    CascadeMux I__3109 (
            .O(N__16918),
            .I(N__16912));
    InMux I__3108 (
            .O(N__16917),
            .I(N__16907));
    InMux I__3107 (
            .O(N__16916),
            .I(N__16907));
    InMux I__3106 (
            .O(N__16915),
            .I(N__16904));
    InMux I__3105 (
            .O(N__16912),
            .I(N__16901));
    LocalMux I__3104 (
            .O(N__16907),
            .I(N__16898));
    LocalMux I__3103 (
            .O(N__16904),
            .I(N__16895));
    LocalMux I__3102 (
            .O(N__16901),
            .I(\sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11 ));
    Odrv4 I__3101 (
            .O(N__16898),
            .I(\sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11 ));
    Odrv4 I__3100 (
            .O(N__16895),
            .I(\sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11 ));
    InMux I__3099 (
            .O(N__16888),
            .I(N__16885));
    LocalMux I__3098 (
            .O(N__16885),
            .I(N__16882));
    Span4Mux_v I__3097 (
            .O(N__16882),
            .I(N__16878));
    InMux I__3096 (
            .O(N__16881),
            .I(N__16875));
    Span4Mux_h I__3095 (
            .O(N__16878),
            .I(N__16872));
    LocalMux I__3094 (
            .O(N__16875),
            .I(\sb_translator_1.cnt19_cry_18_THRU_CO ));
    Odrv4 I__3093 (
            .O(N__16872),
            .I(\sb_translator_1.cnt19_cry_18_THRU_CO ));
    CascadeMux I__3092 (
            .O(N__16867),
            .I(\sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_ ));
    InMux I__3091 (
            .O(N__16864),
            .I(N__16857));
    InMux I__3090 (
            .O(N__16863),
            .I(N__16854));
    InMux I__3089 (
            .O(N__16862),
            .I(N__16845));
    InMux I__3088 (
            .O(N__16861),
            .I(N__16845));
    InMux I__3087 (
            .O(N__16860),
            .I(N__16845));
    LocalMux I__3086 (
            .O(N__16857),
            .I(N__16837));
    LocalMux I__3085 (
            .O(N__16854),
            .I(N__16837));
    InMux I__3084 (
            .O(N__16853),
            .I(N__16834));
    InMux I__3083 (
            .O(N__16852),
            .I(N__16831));
    LocalMux I__3082 (
            .O(N__16845),
            .I(N__16828));
    InMux I__3081 (
            .O(N__16844),
            .I(N__16818));
    InMux I__3080 (
            .O(N__16843),
            .I(N__16818));
    InMux I__3079 (
            .O(N__16842),
            .I(N__16818));
    Span12Mux_h I__3078 (
            .O(N__16837),
            .I(N__16815));
    LocalMux I__3077 (
            .O(N__16834),
            .I(N__16812));
    LocalMux I__3076 (
            .O(N__16831),
            .I(N__16807));
    Span4Mux_h I__3075 (
            .O(N__16828),
            .I(N__16807));
    InMux I__3074 (
            .O(N__16827),
            .I(N__16800));
    InMux I__3073 (
            .O(N__16826),
            .I(N__16800));
    InMux I__3072 (
            .O(N__16825),
            .I(N__16800));
    LocalMux I__3071 (
            .O(N__16818),
            .I(mosi_rx));
    Odrv12 I__3070 (
            .O(N__16815),
            .I(mosi_rx));
    Odrv4 I__3069 (
            .O(N__16812),
            .I(mosi_rx));
    Odrv4 I__3068 (
            .O(N__16807),
            .I(mosi_rx));
    LocalMux I__3067 (
            .O(N__16800),
            .I(mosi_rx));
    CEMux I__3066 (
            .O(N__16789),
            .I(N__16786));
    LocalMux I__3065 (
            .O(N__16786),
            .I(N__16781));
    CEMux I__3064 (
            .O(N__16785),
            .I(N__16778));
    CEMux I__3063 (
            .O(N__16784),
            .I(N__16775));
    Span4Mux_h I__3062 (
            .O(N__16781),
            .I(N__16772));
    LocalMux I__3061 (
            .O(N__16778),
            .I(N__16769));
    LocalMux I__3060 (
            .O(N__16775),
            .I(N__16766));
    Odrv4 I__3059 (
            .O(N__16772),
            .I(\sb_translator_1.state_RNIOH7V9Z0Z_0 ));
    Odrv4 I__3058 (
            .O(N__16769),
            .I(\sb_translator_1.state_RNIOH7V9Z0Z_0 ));
    Odrv4 I__3057 (
            .O(N__16766),
            .I(\sb_translator_1.state_RNIOH7V9Z0Z_0 ));
    InMux I__3056 (
            .O(N__16759),
            .I(N__16756));
    LocalMux I__3055 (
            .O(N__16756),
            .I(N__16753));
    Odrv12 I__3054 (
            .O(N__16753),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_5 ));
    CascadeMux I__3053 (
            .O(N__16750),
            .I(N__16747));
    CascadeBuf I__3052 (
            .O(N__16747),
            .I(N__16744));
    CascadeMux I__3051 (
            .O(N__16744),
            .I(N__16739));
    CascadeMux I__3050 (
            .O(N__16743),
            .I(N__16736));
    CascadeMux I__3049 (
            .O(N__16742),
            .I(N__16733));
    CascadeBuf I__3048 (
            .O(N__16739),
            .I(N__16730));
    CascadeBuf I__3047 (
            .O(N__16736),
            .I(N__16727));
    CascadeBuf I__3046 (
            .O(N__16733),
            .I(N__16723));
    CascadeMux I__3045 (
            .O(N__16730),
            .I(N__16720));
    CascadeMux I__3044 (
            .O(N__16727),
            .I(N__16717));
    CascadeMux I__3043 (
            .O(N__16726),
            .I(N__16714));
    CascadeMux I__3042 (
            .O(N__16723),
            .I(N__16711));
    CascadeBuf I__3041 (
            .O(N__16720),
            .I(N__16708));
    CascadeBuf I__3040 (
            .O(N__16717),
            .I(N__16705));
    CascadeBuf I__3039 (
            .O(N__16714),
            .I(N__16702));
    CascadeBuf I__3038 (
            .O(N__16711),
            .I(N__16699));
    CascadeMux I__3037 (
            .O(N__16708),
            .I(N__16696));
    CascadeMux I__3036 (
            .O(N__16705),
            .I(N__16693));
    CascadeMux I__3035 (
            .O(N__16702),
            .I(N__16690));
    CascadeMux I__3034 (
            .O(N__16699),
            .I(N__16687));
    CascadeBuf I__3033 (
            .O(N__16696),
            .I(N__16684));
    CascadeBuf I__3032 (
            .O(N__16693),
            .I(N__16681));
    CascadeBuf I__3031 (
            .O(N__16690),
            .I(N__16678));
    CascadeBuf I__3030 (
            .O(N__16687),
            .I(N__16675));
    CascadeMux I__3029 (
            .O(N__16684),
            .I(N__16672));
    CascadeMux I__3028 (
            .O(N__16681),
            .I(N__16669));
    CascadeMux I__3027 (
            .O(N__16678),
            .I(N__16666));
    CascadeMux I__3026 (
            .O(N__16675),
            .I(N__16663));
    CascadeBuf I__3025 (
            .O(N__16672),
            .I(N__16660));
    CascadeBuf I__3024 (
            .O(N__16669),
            .I(N__16657));
    CascadeBuf I__3023 (
            .O(N__16666),
            .I(N__16654));
    CascadeBuf I__3022 (
            .O(N__16663),
            .I(N__16651));
    CascadeMux I__3021 (
            .O(N__16660),
            .I(N__16648));
    CascadeMux I__3020 (
            .O(N__16657),
            .I(N__16645));
    CascadeMux I__3019 (
            .O(N__16654),
            .I(N__16642));
    CascadeMux I__3018 (
            .O(N__16651),
            .I(N__16639));
    CascadeBuf I__3017 (
            .O(N__16648),
            .I(N__16636));
    CascadeBuf I__3016 (
            .O(N__16645),
            .I(N__16633));
    CascadeBuf I__3015 (
            .O(N__16642),
            .I(N__16630));
    CascadeBuf I__3014 (
            .O(N__16639),
            .I(N__16627));
    CascadeMux I__3013 (
            .O(N__16636),
            .I(N__16624));
    CascadeMux I__3012 (
            .O(N__16633),
            .I(N__16621));
    CascadeMux I__3011 (
            .O(N__16630),
            .I(N__16618));
    CascadeMux I__3010 (
            .O(N__16627),
            .I(N__16615));
    InMux I__3009 (
            .O(N__16624),
            .I(N__16612));
    CascadeBuf I__3008 (
            .O(N__16621),
            .I(N__16609));
    CascadeBuf I__3007 (
            .O(N__16618),
            .I(N__16606));
    CascadeBuf I__3006 (
            .O(N__16615),
            .I(N__16603));
    LocalMux I__3005 (
            .O(N__16612),
            .I(N__16600));
    CascadeMux I__3004 (
            .O(N__16609),
            .I(N__16597));
    CascadeMux I__3003 (
            .O(N__16606),
            .I(N__16594));
    CascadeMux I__3002 (
            .O(N__16603),
            .I(N__16591));
    Span4Mux_s1_v I__3001 (
            .O(N__16600),
            .I(N__16587));
    InMux I__3000 (
            .O(N__16597),
            .I(N__16584));
    CascadeBuf I__2999 (
            .O(N__16594),
            .I(N__16581));
    InMux I__2998 (
            .O(N__16591),
            .I(N__16578));
    InMux I__2997 (
            .O(N__16590),
            .I(N__16575));
    Span4Mux_s2_h I__2996 (
            .O(N__16587),
            .I(N__16570));
    LocalMux I__2995 (
            .O(N__16584),
            .I(N__16570));
    CascadeMux I__2994 (
            .O(N__16581),
            .I(N__16567));
    LocalMux I__2993 (
            .O(N__16578),
            .I(N__16564));
    LocalMux I__2992 (
            .O(N__16575),
            .I(N__16559));
    Span4Mux_h I__2991 (
            .O(N__16570),
            .I(N__16559));
    InMux I__2990 (
            .O(N__16567),
            .I(N__16556));
    Span4Mux_s1_v I__2989 (
            .O(N__16564),
            .I(N__16549));
    Span4Mux_h I__2988 (
            .O(N__16559),
            .I(N__16549));
    LocalMux I__2987 (
            .O(N__16556),
            .I(N__16549));
    Span4Mux_v I__2986 (
            .O(N__16549),
            .I(N__16546));
    Span4Mux_v I__2985 (
            .O(N__16546),
            .I(N__16543));
    Odrv4 I__2984 (
            .O(N__16543),
            .I(addr_out_5));
    CascadeMux I__2983 (
            .O(N__16540),
            .I(N__16535));
    CascadeMux I__2982 (
            .O(N__16539),
            .I(N__16532));
    CascadeMux I__2981 (
            .O(N__16538),
            .I(N__16529));
    CascadeBuf I__2980 (
            .O(N__16535),
            .I(N__16526));
    CascadeBuf I__2979 (
            .O(N__16532),
            .I(N__16522));
    CascadeBuf I__2978 (
            .O(N__16529),
            .I(N__16519));
    CascadeMux I__2977 (
            .O(N__16526),
            .I(N__16516));
    CascadeMux I__2976 (
            .O(N__16525),
            .I(N__16513));
    CascadeMux I__2975 (
            .O(N__16522),
            .I(N__16510));
    CascadeMux I__2974 (
            .O(N__16519),
            .I(N__16507));
    CascadeBuf I__2973 (
            .O(N__16516),
            .I(N__16504));
    CascadeBuf I__2972 (
            .O(N__16513),
            .I(N__16501));
    CascadeBuf I__2971 (
            .O(N__16510),
            .I(N__16498));
    CascadeBuf I__2970 (
            .O(N__16507),
            .I(N__16495));
    CascadeMux I__2969 (
            .O(N__16504),
            .I(N__16492));
    CascadeMux I__2968 (
            .O(N__16501),
            .I(N__16489));
    CascadeMux I__2967 (
            .O(N__16498),
            .I(N__16486));
    CascadeMux I__2966 (
            .O(N__16495),
            .I(N__16483));
    CascadeBuf I__2965 (
            .O(N__16492),
            .I(N__16480));
    CascadeBuf I__2964 (
            .O(N__16489),
            .I(N__16477));
    CascadeBuf I__2963 (
            .O(N__16486),
            .I(N__16474));
    CascadeBuf I__2962 (
            .O(N__16483),
            .I(N__16471));
    CascadeMux I__2961 (
            .O(N__16480),
            .I(N__16468));
    CascadeMux I__2960 (
            .O(N__16477),
            .I(N__16465));
    CascadeMux I__2959 (
            .O(N__16474),
            .I(N__16462));
    CascadeMux I__2958 (
            .O(N__16471),
            .I(N__16459));
    CascadeBuf I__2957 (
            .O(N__16468),
            .I(N__16456));
    CascadeBuf I__2956 (
            .O(N__16465),
            .I(N__16453));
    CascadeBuf I__2955 (
            .O(N__16462),
            .I(N__16450));
    CascadeBuf I__2954 (
            .O(N__16459),
            .I(N__16447));
    CascadeMux I__2953 (
            .O(N__16456),
            .I(N__16444));
    CascadeMux I__2952 (
            .O(N__16453),
            .I(N__16441));
    CascadeMux I__2951 (
            .O(N__16450),
            .I(N__16438));
    CascadeMux I__2950 (
            .O(N__16447),
            .I(N__16435));
    CascadeBuf I__2949 (
            .O(N__16444),
            .I(N__16432));
    CascadeBuf I__2948 (
            .O(N__16441),
            .I(N__16429));
    CascadeBuf I__2947 (
            .O(N__16438),
            .I(N__16426));
    CascadeBuf I__2946 (
            .O(N__16435),
            .I(N__16423));
    CascadeMux I__2945 (
            .O(N__16432),
            .I(N__16420));
    CascadeMux I__2944 (
            .O(N__16429),
            .I(N__16417));
    CascadeMux I__2943 (
            .O(N__16426),
            .I(N__16414));
    CascadeMux I__2942 (
            .O(N__16423),
            .I(N__16411));
    CascadeBuf I__2941 (
            .O(N__16420),
            .I(N__16408));
    CascadeBuf I__2940 (
            .O(N__16417),
            .I(N__16405));
    CascadeBuf I__2939 (
            .O(N__16414),
            .I(N__16402));
    CascadeBuf I__2938 (
            .O(N__16411),
            .I(N__16399));
    CascadeMux I__2937 (
            .O(N__16408),
            .I(N__16396));
    CascadeMux I__2936 (
            .O(N__16405),
            .I(N__16393));
    CascadeMux I__2935 (
            .O(N__16402),
            .I(N__16390));
    CascadeMux I__2934 (
            .O(N__16399),
            .I(N__16387));
    InMux I__2933 (
            .O(N__16396),
            .I(N__16383));
    CascadeBuf I__2932 (
            .O(N__16393),
            .I(N__16380));
    InMux I__2931 (
            .O(N__16390),
            .I(N__16377));
    InMux I__2930 (
            .O(N__16387),
            .I(N__16374));
    InMux I__2929 (
            .O(N__16386),
            .I(N__16371));
    LocalMux I__2928 (
            .O(N__16383),
            .I(N__16368));
    CascadeMux I__2927 (
            .O(N__16380),
            .I(N__16365));
    LocalMux I__2926 (
            .O(N__16377),
            .I(N__16362));
    LocalMux I__2925 (
            .O(N__16374),
            .I(N__16359));
    LocalMux I__2924 (
            .O(N__16371),
            .I(N__16354));
    Span4Mux_h I__2923 (
            .O(N__16368),
            .I(N__16354));
    InMux I__2922 (
            .O(N__16365),
            .I(N__16351));
    Span4Mux_s3_v I__2921 (
            .O(N__16362),
            .I(N__16348));
    Span4Mux_s1_v I__2920 (
            .O(N__16359),
            .I(N__16341));
    Span4Mux_h I__2919 (
            .O(N__16354),
            .I(N__16341));
    LocalMux I__2918 (
            .O(N__16351),
            .I(N__16341));
    Span4Mux_v I__2917 (
            .O(N__16348),
            .I(N__16338));
    Span4Mux_v I__2916 (
            .O(N__16341),
            .I(N__16335));
    Span4Mux_h I__2915 (
            .O(N__16338),
            .I(N__16332));
    Span4Mux_v I__2914 (
            .O(N__16335),
            .I(N__16329));
    Odrv4 I__2913 (
            .O(N__16332),
            .I(addr_out_6));
    Odrv4 I__2912 (
            .O(N__16329),
            .I(addr_out_6));
    CascadeMux I__2911 (
            .O(N__16324),
            .I(N__16319));
    CascadeMux I__2910 (
            .O(N__16323),
            .I(N__16316));
    CascadeMux I__2909 (
            .O(N__16322),
            .I(N__16313));
    CascadeBuf I__2908 (
            .O(N__16319),
            .I(N__16310));
    CascadeBuf I__2907 (
            .O(N__16316),
            .I(N__16306));
    CascadeBuf I__2906 (
            .O(N__16313),
            .I(N__16303));
    CascadeMux I__2905 (
            .O(N__16310),
            .I(N__16300));
    CascadeMux I__2904 (
            .O(N__16309),
            .I(N__16297));
    CascadeMux I__2903 (
            .O(N__16306),
            .I(N__16294));
    CascadeMux I__2902 (
            .O(N__16303),
            .I(N__16291));
    CascadeBuf I__2901 (
            .O(N__16300),
            .I(N__16288));
    CascadeBuf I__2900 (
            .O(N__16297),
            .I(N__16285));
    CascadeBuf I__2899 (
            .O(N__16294),
            .I(N__16282));
    CascadeBuf I__2898 (
            .O(N__16291),
            .I(N__16279));
    CascadeMux I__2897 (
            .O(N__16288),
            .I(N__16276));
    CascadeMux I__2896 (
            .O(N__16285),
            .I(N__16273));
    CascadeMux I__2895 (
            .O(N__16282),
            .I(N__16270));
    CascadeMux I__2894 (
            .O(N__16279),
            .I(N__16267));
    CascadeBuf I__2893 (
            .O(N__16276),
            .I(N__16264));
    CascadeBuf I__2892 (
            .O(N__16273),
            .I(N__16261));
    CascadeBuf I__2891 (
            .O(N__16270),
            .I(N__16258));
    CascadeBuf I__2890 (
            .O(N__16267),
            .I(N__16255));
    CascadeMux I__2889 (
            .O(N__16264),
            .I(N__16252));
    CascadeMux I__2888 (
            .O(N__16261),
            .I(N__16249));
    CascadeMux I__2887 (
            .O(N__16258),
            .I(N__16246));
    CascadeMux I__2886 (
            .O(N__16255),
            .I(N__16243));
    CascadeBuf I__2885 (
            .O(N__16252),
            .I(N__16240));
    CascadeBuf I__2884 (
            .O(N__16249),
            .I(N__16237));
    CascadeBuf I__2883 (
            .O(N__16246),
            .I(N__16234));
    CascadeBuf I__2882 (
            .O(N__16243),
            .I(N__16231));
    CascadeMux I__2881 (
            .O(N__16240),
            .I(N__16228));
    CascadeMux I__2880 (
            .O(N__16237),
            .I(N__16225));
    CascadeMux I__2879 (
            .O(N__16234),
            .I(N__16222));
    CascadeMux I__2878 (
            .O(N__16231),
            .I(N__16219));
    CascadeBuf I__2877 (
            .O(N__16228),
            .I(N__16216));
    CascadeBuf I__2876 (
            .O(N__16225),
            .I(N__16213));
    CascadeBuf I__2875 (
            .O(N__16222),
            .I(N__16210));
    CascadeBuf I__2874 (
            .O(N__16219),
            .I(N__16207));
    CascadeMux I__2873 (
            .O(N__16216),
            .I(N__16204));
    CascadeMux I__2872 (
            .O(N__16213),
            .I(N__16201));
    CascadeMux I__2871 (
            .O(N__16210),
            .I(N__16198));
    CascadeMux I__2870 (
            .O(N__16207),
            .I(N__16195));
    CascadeBuf I__2869 (
            .O(N__16204),
            .I(N__16192));
    CascadeBuf I__2868 (
            .O(N__16201),
            .I(N__16189));
    CascadeBuf I__2867 (
            .O(N__16198),
            .I(N__16186));
    CascadeBuf I__2866 (
            .O(N__16195),
            .I(N__16183));
    CascadeMux I__2865 (
            .O(N__16192),
            .I(N__16180));
    CascadeMux I__2864 (
            .O(N__16189),
            .I(N__16177));
    CascadeMux I__2863 (
            .O(N__16186),
            .I(N__16174));
    CascadeMux I__2862 (
            .O(N__16183),
            .I(N__16171));
    InMux I__2861 (
            .O(N__16180),
            .I(N__16167));
    CascadeBuf I__2860 (
            .O(N__16177),
            .I(N__16164));
    InMux I__2859 (
            .O(N__16174),
            .I(N__16161));
    InMux I__2858 (
            .O(N__16171),
            .I(N__16158));
    InMux I__2857 (
            .O(N__16170),
            .I(N__16155));
    LocalMux I__2856 (
            .O(N__16167),
            .I(N__16152));
    CascadeMux I__2855 (
            .O(N__16164),
            .I(N__16149));
    LocalMux I__2854 (
            .O(N__16161),
            .I(N__16146));
    LocalMux I__2853 (
            .O(N__16158),
            .I(N__16143));
    LocalMux I__2852 (
            .O(N__16155),
            .I(N__16138));
    Span4Mux_h I__2851 (
            .O(N__16152),
            .I(N__16138));
    InMux I__2850 (
            .O(N__16149),
            .I(N__16135));
    Span4Mux_s2_v I__2849 (
            .O(N__16146),
            .I(N__16132));
    Span4Mux_s1_v I__2848 (
            .O(N__16143),
            .I(N__16125));
    Span4Mux_h I__2847 (
            .O(N__16138),
            .I(N__16125));
    LocalMux I__2846 (
            .O(N__16135),
            .I(N__16125));
    Span4Mux_h I__2845 (
            .O(N__16132),
            .I(N__16122));
    Span4Mux_v I__2844 (
            .O(N__16125),
            .I(N__16119));
    Span4Mux_v I__2843 (
            .O(N__16122),
            .I(N__16116));
    Span4Mux_v I__2842 (
            .O(N__16119),
            .I(N__16113));
    Odrv4 I__2841 (
            .O(N__16116),
            .I(addr_out_7));
    Odrv4 I__2840 (
            .O(N__16113),
            .I(addr_out_7));
    InMux I__2839 (
            .O(N__16108),
            .I(N__16105));
    LocalMux I__2838 (
            .O(N__16105),
            .I(N__16100));
    CascadeMux I__2837 (
            .O(N__16104),
            .I(N__16096));
    CascadeMux I__2836 (
            .O(N__16103),
            .I(N__16093));
    Span4Mux_h I__2835 (
            .O(N__16100),
            .I(N__16090));
    InMux I__2834 (
            .O(N__16099),
            .I(N__16083));
    InMux I__2833 (
            .O(N__16096),
            .I(N__16083));
    InMux I__2832 (
            .O(N__16093),
            .I(N__16083));
    Odrv4 I__2831 (
            .O(N__16090),
            .I(\sb_translator_1.cnt_RNILAHE_2Z0Z_10 ));
    LocalMux I__2830 (
            .O(N__16083),
            .I(\sb_translator_1.cnt_RNILAHE_2Z0Z_10 ));
    InMux I__2829 (
            .O(N__16078),
            .I(N__16072));
    InMux I__2828 (
            .O(N__16077),
            .I(N__16072));
    LocalMux I__2827 (
            .O(N__16072),
            .I(N__16067));
    InMux I__2826 (
            .O(N__16071),
            .I(N__16062));
    InMux I__2825 (
            .O(N__16070),
            .I(N__16062));
    Span4Mux_v I__2824 (
            .O(N__16067),
            .I(N__16057));
    LocalMux I__2823 (
            .O(N__16062),
            .I(N__16057));
    Odrv4 I__2822 (
            .O(N__16057),
            .I(\sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10 ));
    CascadeMux I__2821 (
            .O(N__16054),
            .I(N__16050));
    CascadeMux I__2820 (
            .O(N__16053),
            .I(N__16046));
    InMux I__2819 (
            .O(N__16050),
            .I(N__16039));
    InMux I__2818 (
            .O(N__16049),
            .I(N__16039));
    InMux I__2817 (
            .O(N__16046),
            .I(N__16039));
    LocalMux I__2816 (
            .O(N__16039),
            .I(N__16035));
    InMux I__2815 (
            .O(N__16038),
            .I(N__16032));
    Span4Mux_v I__2814 (
            .O(N__16035),
            .I(N__16027));
    LocalMux I__2813 (
            .O(N__16032),
            .I(N__16027));
    Odrv4 I__2812 (
            .O(N__16027),
            .I(\sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10 ));
    InMux I__2811 (
            .O(N__16024),
            .I(N__16019));
    InMux I__2810 (
            .O(N__16023),
            .I(N__16016));
    InMux I__2809 (
            .O(N__16022),
            .I(N__16013));
    LocalMux I__2808 (
            .O(N__16019),
            .I(N__16010));
    LocalMux I__2807 (
            .O(N__16016),
            .I(mosi_data_out_0));
    LocalMux I__2806 (
            .O(N__16013),
            .I(mosi_data_out_0));
    Odrv4 I__2805 (
            .O(N__16010),
            .I(mosi_data_out_0));
    InMux I__2804 (
            .O(N__16003),
            .I(N__16000));
    LocalMux I__2803 (
            .O(N__16000),
            .I(\sb_translator_1.instr_tmpZ1Z_0 ));
    InMux I__2802 (
            .O(N__15997),
            .I(N__15993));
    InMux I__2801 (
            .O(N__15996),
            .I(N__15990));
    LocalMux I__2800 (
            .O(N__15993),
            .I(N__15986));
    LocalMux I__2799 (
            .O(N__15990),
            .I(N__15983));
    InMux I__2798 (
            .O(N__15989),
            .I(N__15980));
    Span4Mux_v I__2797 (
            .O(N__15986),
            .I(N__15973));
    Span4Mux_h I__2796 (
            .O(N__15983),
            .I(N__15973));
    LocalMux I__2795 (
            .O(N__15980),
            .I(N__15973));
    Span4Mux_h I__2794 (
            .O(N__15973),
            .I(N__15970));
    Odrv4 I__2793 (
            .O(N__15970),
            .I(mosi_data_out_1));
    InMux I__2792 (
            .O(N__15967),
            .I(N__15964));
    LocalMux I__2791 (
            .O(N__15964),
            .I(\sb_translator_1.instr_tmpZ1Z_1 ));
    InMux I__2790 (
            .O(N__15961),
            .I(N__15958));
    LocalMux I__2789 (
            .O(N__15958),
            .I(N__15953));
    InMux I__2788 (
            .O(N__15957),
            .I(N__15950));
    InMux I__2787 (
            .O(N__15956),
            .I(N__15947));
    Odrv4 I__2786 (
            .O(N__15953),
            .I(mosi_data_out_2));
    LocalMux I__2785 (
            .O(N__15950),
            .I(mosi_data_out_2));
    LocalMux I__2784 (
            .O(N__15947),
            .I(mosi_data_out_2));
    InMux I__2783 (
            .O(N__15940),
            .I(N__15937));
    LocalMux I__2782 (
            .O(N__15937),
            .I(\sb_translator_1.instr_tmpZ1Z_2 ));
    CascadeMux I__2781 (
            .O(N__15934),
            .I(N__15929));
    CascadeMux I__2780 (
            .O(N__15933),
            .I(N__15925));
    InMux I__2779 (
            .O(N__15932),
            .I(N__15918));
    InMux I__2778 (
            .O(N__15929),
            .I(N__15918));
    InMux I__2777 (
            .O(N__15928),
            .I(N__15913));
    InMux I__2776 (
            .O(N__15925),
            .I(N__15913));
    InMux I__2775 (
            .O(N__15924),
            .I(N__15908));
    InMux I__2774 (
            .O(N__15923),
            .I(N__15908));
    LocalMux I__2773 (
            .O(N__15918),
            .I(\sb_translator_1.num_ledsZ0Z_9 ));
    LocalMux I__2772 (
            .O(N__15913),
            .I(\sb_translator_1.num_ledsZ0Z_9 ));
    LocalMux I__2771 (
            .O(N__15908),
            .I(\sb_translator_1.num_ledsZ0Z_9 ));
    CascadeMux I__2770 (
            .O(N__15901),
            .I(N__15897));
    InMux I__2769 (
            .O(N__15900),
            .I(N__15888));
    InMux I__2768 (
            .O(N__15897),
            .I(N__15888));
    InMux I__2767 (
            .O(N__15896),
            .I(N__15879));
    InMux I__2766 (
            .O(N__15895),
            .I(N__15879));
    InMux I__2765 (
            .O(N__15894),
            .I(N__15879));
    InMux I__2764 (
            .O(N__15893),
            .I(N__15879));
    LocalMux I__2763 (
            .O(N__15888),
            .I(\sb_translator_1.num_ledsZ0Z_11 ));
    LocalMux I__2762 (
            .O(N__15879),
            .I(\sb_translator_1.num_ledsZ0Z_11 ));
    CascadeMux I__2761 (
            .O(N__15874),
            .I(N__15869));
    CascadeMux I__2760 (
            .O(N__15873),
            .I(N__15864));
    InMux I__2759 (
            .O(N__15872),
            .I(N__15858));
    InMux I__2758 (
            .O(N__15869),
            .I(N__15858));
    InMux I__2757 (
            .O(N__15868),
            .I(N__15849));
    InMux I__2756 (
            .O(N__15867),
            .I(N__15849));
    InMux I__2755 (
            .O(N__15864),
            .I(N__15849));
    InMux I__2754 (
            .O(N__15863),
            .I(N__15849));
    LocalMux I__2753 (
            .O(N__15858),
            .I(\sb_translator_1.num_ledsZ0Z_10 ));
    LocalMux I__2752 (
            .O(N__15849),
            .I(\sb_translator_1.num_ledsZ0Z_10 ));
    CascadeMux I__2751 (
            .O(N__15844),
            .I(\sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_ ));
    InMux I__2750 (
            .O(N__15841),
            .I(N__15837));
    InMux I__2749 (
            .O(N__15840),
            .I(N__15834));
    LocalMux I__2748 (
            .O(N__15837),
            .I(N__15831));
    LocalMux I__2747 (
            .O(N__15834),
            .I(N__15828));
    Span4Mux_v I__2746 (
            .O(N__15831),
            .I(N__15823));
    Span4Mux_v I__2745 (
            .O(N__15828),
            .I(N__15823));
    Odrv4 I__2744 (
            .O(N__15823),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_0_0_7 ));
    InMux I__2743 (
            .O(N__15820),
            .I(N__15815));
    InMux I__2742 (
            .O(N__15819),
            .I(N__15810));
    InMux I__2741 (
            .O(N__15818),
            .I(N__15810));
    LocalMux I__2740 (
            .O(N__15815),
            .I(N__15804));
    LocalMux I__2739 (
            .O(N__15810),
            .I(N__15804));
    InMux I__2738 (
            .O(N__15809),
            .I(N__15801));
    Span4Mux_v I__2737 (
            .O(N__15804),
            .I(N__15796));
    LocalMux I__2736 (
            .O(N__15801),
            .I(N__15796));
    Span4Mux_v I__2735 (
            .O(N__15796),
            .I(N__15793));
    Odrv4 I__2734 (
            .O(N__15793),
            .I(\sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10 ));
    InMux I__2733 (
            .O(N__15790),
            .I(N__15787));
    LocalMux I__2732 (
            .O(N__15787),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_0 ));
    CascadeMux I__2731 (
            .O(N__15784),
            .I(N__15781));
    CascadeBuf I__2730 (
            .O(N__15781),
            .I(N__15777));
    CascadeMux I__2729 (
            .O(N__15780),
            .I(N__15774));
    CascadeMux I__2728 (
            .O(N__15777),
            .I(N__15770));
    CascadeBuf I__2727 (
            .O(N__15774),
            .I(N__15767));
    CascadeMux I__2726 (
            .O(N__15773),
            .I(N__15763));
    CascadeBuf I__2725 (
            .O(N__15770),
            .I(N__15760));
    CascadeMux I__2724 (
            .O(N__15767),
            .I(N__15757));
    CascadeMux I__2723 (
            .O(N__15766),
            .I(N__15754));
    CascadeBuf I__2722 (
            .O(N__15763),
            .I(N__15751));
    CascadeMux I__2721 (
            .O(N__15760),
            .I(N__15748));
    CascadeBuf I__2720 (
            .O(N__15757),
            .I(N__15745));
    CascadeBuf I__2719 (
            .O(N__15754),
            .I(N__15742));
    CascadeMux I__2718 (
            .O(N__15751),
            .I(N__15739));
    CascadeBuf I__2717 (
            .O(N__15748),
            .I(N__15736));
    CascadeMux I__2716 (
            .O(N__15745),
            .I(N__15733));
    CascadeMux I__2715 (
            .O(N__15742),
            .I(N__15730));
    CascadeBuf I__2714 (
            .O(N__15739),
            .I(N__15727));
    CascadeMux I__2713 (
            .O(N__15736),
            .I(N__15724));
    CascadeBuf I__2712 (
            .O(N__15733),
            .I(N__15721));
    CascadeBuf I__2711 (
            .O(N__15730),
            .I(N__15718));
    CascadeMux I__2710 (
            .O(N__15727),
            .I(N__15715));
    CascadeBuf I__2709 (
            .O(N__15724),
            .I(N__15712));
    CascadeMux I__2708 (
            .O(N__15721),
            .I(N__15709));
    CascadeMux I__2707 (
            .O(N__15718),
            .I(N__15706));
    CascadeBuf I__2706 (
            .O(N__15715),
            .I(N__15703));
    CascadeMux I__2705 (
            .O(N__15712),
            .I(N__15700));
    CascadeBuf I__2704 (
            .O(N__15709),
            .I(N__15697));
    CascadeBuf I__2703 (
            .O(N__15706),
            .I(N__15694));
    CascadeMux I__2702 (
            .O(N__15703),
            .I(N__15691));
    CascadeBuf I__2701 (
            .O(N__15700),
            .I(N__15688));
    CascadeMux I__2700 (
            .O(N__15697),
            .I(N__15685));
    CascadeMux I__2699 (
            .O(N__15694),
            .I(N__15682));
    CascadeBuf I__2698 (
            .O(N__15691),
            .I(N__15679));
    CascadeMux I__2697 (
            .O(N__15688),
            .I(N__15676));
    CascadeBuf I__2696 (
            .O(N__15685),
            .I(N__15673));
    CascadeBuf I__2695 (
            .O(N__15682),
            .I(N__15670));
    CascadeMux I__2694 (
            .O(N__15679),
            .I(N__15667));
    CascadeBuf I__2693 (
            .O(N__15676),
            .I(N__15664));
    CascadeMux I__2692 (
            .O(N__15673),
            .I(N__15661));
    CascadeMux I__2691 (
            .O(N__15670),
            .I(N__15658));
    CascadeBuf I__2690 (
            .O(N__15667),
            .I(N__15655));
    CascadeMux I__2689 (
            .O(N__15664),
            .I(N__15652));
    CascadeBuf I__2688 (
            .O(N__15661),
            .I(N__15649));
    CascadeBuf I__2687 (
            .O(N__15658),
            .I(N__15646));
    CascadeMux I__2686 (
            .O(N__15655),
            .I(N__15643));
    InMux I__2685 (
            .O(N__15652),
            .I(N__15640));
    CascadeMux I__2684 (
            .O(N__15649),
            .I(N__15637));
    CascadeMux I__2683 (
            .O(N__15646),
            .I(N__15634));
    CascadeBuf I__2682 (
            .O(N__15643),
            .I(N__15631));
    LocalMux I__2681 (
            .O(N__15640),
            .I(N__15628));
    InMux I__2680 (
            .O(N__15637),
            .I(N__15625));
    CascadeBuf I__2679 (
            .O(N__15634),
            .I(N__15622));
    CascadeMux I__2678 (
            .O(N__15631),
            .I(N__15618));
    Span4Mux_s1_v I__2677 (
            .O(N__15628),
            .I(N__15615));
    LocalMux I__2676 (
            .O(N__15625),
            .I(N__15612));
    CascadeMux I__2675 (
            .O(N__15622),
            .I(N__15609));
    InMux I__2674 (
            .O(N__15621),
            .I(N__15606));
    InMux I__2673 (
            .O(N__15618),
            .I(N__15603));
    Span4Mux_h I__2672 (
            .O(N__15615),
            .I(N__15598));
    Span4Mux_s1_v I__2671 (
            .O(N__15612),
            .I(N__15598));
    InMux I__2670 (
            .O(N__15609),
            .I(N__15595));
    LocalMux I__2669 (
            .O(N__15606),
            .I(N__15592));
    LocalMux I__2668 (
            .O(N__15603),
            .I(N__15589));
    Sp12to4 I__2667 (
            .O(N__15598),
            .I(N__15584));
    LocalMux I__2666 (
            .O(N__15595),
            .I(N__15584));
    Span12Mux_s9_v I__2665 (
            .O(N__15592),
            .I(N__15581));
    Span12Mux_s7_h I__2664 (
            .O(N__15589),
            .I(N__15576));
    Span12Mux_s6_h I__2663 (
            .O(N__15584),
            .I(N__15576));
    Odrv12 I__2662 (
            .O(N__15581),
            .I(addr_out_0));
    Odrv12 I__2661 (
            .O(N__15576),
            .I(addr_out_0));
    CascadeMux I__2660 (
            .O(N__15571),
            .I(N__15568));
    InMux I__2659 (
            .O(N__15568),
            .I(N__15565));
    LocalMux I__2658 (
            .O(N__15565),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_1 ));
    CascadeMux I__2657 (
            .O(N__15562),
            .I(N__15558));
    CascadeMux I__2656 (
            .O(N__15561),
            .I(N__15555));
    CascadeBuf I__2655 (
            .O(N__15558),
            .I(N__15550));
    CascadeBuf I__2654 (
            .O(N__15555),
            .I(N__15547));
    CascadeMux I__2653 (
            .O(N__15554),
            .I(N__15544));
    CascadeMux I__2652 (
            .O(N__15553),
            .I(N__15541));
    CascadeMux I__2651 (
            .O(N__15550),
            .I(N__15538));
    CascadeMux I__2650 (
            .O(N__15547),
            .I(N__15535));
    CascadeBuf I__2649 (
            .O(N__15544),
            .I(N__15532));
    CascadeBuf I__2648 (
            .O(N__15541),
            .I(N__15529));
    CascadeBuf I__2647 (
            .O(N__15538),
            .I(N__15526));
    CascadeBuf I__2646 (
            .O(N__15535),
            .I(N__15523));
    CascadeMux I__2645 (
            .O(N__15532),
            .I(N__15520));
    CascadeMux I__2644 (
            .O(N__15529),
            .I(N__15517));
    CascadeMux I__2643 (
            .O(N__15526),
            .I(N__15514));
    CascadeMux I__2642 (
            .O(N__15523),
            .I(N__15511));
    CascadeBuf I__2641 (
            .O(N__15520),
            .I(N__15508));
    CascadeBuf I__2640 (
            .O(N__15517),
            .I(N__15505));
    CascadeBuf I__2639 (
            .O(N__15514),
            .I(N__15502));
    CascadeBuf I__2638 (
            .O(N__15511),
            .I(N__15499));
    CascadeMux I__2637 (
            .O(N__15508),
            .I(N__15496));
    CascadeMux I__2636 (
            .O(N__15505),
            .I(N__15493));
    CascadeMux I__2635 (
            .O(N__15502),
            .I(N__15490));
    CascadeMux I__2634 (
            .O(N__15499),
            .I(N__15487));
    CascadeBuf I__2633 (
            .O(N__15496),
            .I(N__15484));
    CascadeBuf I__2632 (
            .O(N__15493),
            .I(N__15481));
    CascadeBuf I__2631 (
            .O(N__15490),
            .I(N__15478));
    CascadeBuf I__2630 (
            .O(N__15487),
            .I(N__15475));
    CascadeMux I__2629 (
            .O(N__15484),
            .I(N__15472));
    CascadeMux I__2628 (
            .O(N__15481),
            .I(N__15469));
    CascadeMux I__2627 (
            .O(N__15478),
            .I(N__15466));
    CascadeMux I__2626 (
            .O(N__15475),
            .I(N__15463));
    CascadeBuf I__2625 (
            .O(N__15472),
            .I(N__15460));
    CascadeBuf I__2624 (
            .O(N__15469),
            .I(N__15457));
    CascadeBuf I__2623 (
            .O(N__15466),
            .I(N__15454));
    CascadeBuf I__2622 (
            .O(N__15463),
            .I(N__15451));
    CascadeMux I__2621 (
            .O(N__15460),
            .I(N__15448));
    CascadeMux I__2620 (
            .O(N__15457),
            .I(N__15445));
    CascadeMux I__2619 (
            .O(N__15454),
            .I(N__15442));
    CascadeMux I__2618 (
            .O(N__15451),
            .I(N__15439));
    CascadeBuf I__2617 (
            .O(N__15448),
            .I(N__15436));
    CascadeBuf I__2616 (
            .O(N__15445),
            .I(N__15433));
    CascadeBuf I__2615 (
            .O(N__15442),
            .I(N__15430));
    CascadeBuf I__2614 (
            .O(N__15439),
            .I(N__15427));
    CascadeMux I__2613 (
            .O(N__15436),
            .I(N__15424));
    CascadeMux I__2612 (
            .O(N__15433),
            .I(N__15421));
    CascadeMux I__2611 (
            .O(N__15430),
            .I(N__15418));
    CascadeMux I__2610 (
            .O(N__15427),
            .I(N__15415));
    CascadeBuf I__2609 (
            .O(N__15424),
            .I(N__15412));
    CascadeBuf I__2608 (
            .O(N__15421),
            .I(N__15409));
    InMux I__2607 (
            .O(N__15418),
            .I(N__15405));
    InMux I__2606 (
            .O(N__15415),
            .I(N__15402));
    CascadeMux I__2605 (
            .O(N__15412),
            .I(N__15399));
    CascadeMux I__2604 (
            .O(N__15409),
            .I(N__15396));
    InMux I__2603 (
            .O(N__15408),
            .I(N__15393));
    LocalMux I__2602 (
            .O(N__15405),
            .I(N__15388));
    LocalMux I__2601 (
            .O(N__15402),
            .I(N__15388));
    InMux I__2600 (
            .O(N__15399),
            .I(N__15385));
    InMux I__2599 (
            .O(N__15396),
            .I(N__15382));
    LocalMux I__2598 (
            .O(N__15393),
            .I(N__15379));
    Span4Mux_s3_v I__2597 (
            .O(N__15388),
            .I(N__15376));
    LocalMux I__2596 (
            .O(N__15385),
            .I(N__15371));
    LocalMux I__2595 (
            .O(N__15382),
            .I(N__15371));
    Span4Mux_v I__2594 (
            .O(N__15379),
            .I(N__15364));
    Span4Mux_h I__2593 (
            .O(N__15376),
            .I(N__15364));
    Span4Mux_s3_v I__2592 (
            .O(N__15371),
            .I(N__15364));
    Span4Mux_h I__2591 (
            .O(N__15364),
            .I(N__15361));
    Span4Mux_v I__2590 (
            .O(N__15361),
            .I(N__15358));
    Odrv4 I__2589 (
            .O(N__15358),
            .I(addr_out_1));
    InMux I__2588 (
            .O(N__15355),
            .I(N__15352));
    LocalMux I__2587 (
            .O(N__15352),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_2 ));
    CascadeMux I__2586 (
            .O(N__15349),
            .I(N__15346));
    CascadeBuf I__2585 (
            .O(N__15346),
            .I(N__15343));
    CascadeMux I__2584 (
            .O(N__15343),
            .I(N__15338));
    CascadeMux I__2583 (
            .O(N__15342),
            .I(N__15335));
    CascadeMux I__2582 (
            .O(N__15341),
            .I(N__15332));
    CascadeBuf I__2581 (
            .O(N__15338),
            .I(N__15329));
    CascadeBuf I__2580 (
            .O(N__15335),
            .I(N__15326));
    CascadeBuf I__2579 (
            .O(N__15332),
            .I(N__15322));
    CascadeMux I__2578 (
            .O(N__15329),
            .I(N__15319));
    CascadeMux I__2577 (
            .O(N__15326),
            .I(N__15316));
    CascadeMux I__2576 (
            .O(N__15325),
            .I(N__15313));
    CascadeMux I__2575 (
            .O(N__15322),
            .I(N__15310));
    CascadeBuf I__2574 (
            .O(N__15319),
            .I(N__15307));
    CascadeBuf I__2573 (
            .O(N__15316),
            .I(N__15304));
    CascadeBuf I__2572 (
            .O(N__15313),
            .I(N__15301));
    CascadeBuf I__2571 (
            .O(N__15310),
            .I(N__15298));
    CascadeMux I__2570 (
            .O(N__15307),
            .I(N__15295));
    CascadeMux I__2569 (
            .O(N__15304),
            .I(N__15292));
    CascadeMux I__2568 (
            .O(N__15301),
            .I(N__15289));
    CascadeMux I__2567 (
            .O(N__15298),
            .I(N__15286));
    CascadeBuf I__2566 (
            .O(N__15295),
            .I(N__15283));
    CascadeBuf I__2565 (
            .O(N__15292),
            .I(N__15280));
    CascadeBuf I__2564 (
            .O(N__15289),
            .I(N__15277));
    CascadeBuf I__2563 (
            .O(N__15286),
            .I(N__15274));
    CascadeMux I__2562 (
            .O(N__15283),
            .I(N__15271));
    CascadeMux I__2561 (
            .O(N__15280),
            .I(N__15268));
    CascadeMux I__2560 (
            .O(N__15277),
            .I(N__15265));
    CascadeMux I__2559 (
            .O(N__15274),
            .I(N__15262));
    CascadeBuf I__2558 (
            .O(N__15271),
            .I(N__15259));
    CascadeBuf I__2557 (
            .O(N__15268),
            .I(N__15256));
    CascadeBuf I__2556 (
            .O(N__15265),
            .I(N__15253));
    CascadeBuf I__2555 (
            .O(N__15262),
            .I(N__15250));
    CascadeMux I__2554 (
            .O(N__15259),
            .I(N__15247));
    CascadeMux I__2553 (
            .O(N__15256),
            .I(N__15244));
    CascadeMux I__2552 (
            .O(N__15253),
            .I(N__15241));
    CascadeMux I__2551 (
            .O(N__15250),
            .I(N__15238));
    CascadeBuf I__2550 (
            .O(N__15247),
            .I(N__15235));
    CascadeBuf I__2549 (
            .O(N__15244),
            .I(N__15232));
    CascadeBuf I__2548 (
            .O(N__15241),
            .I(N__15229));
    CascadeBuf I__2547 (
            .O(N__15238),
            .I(N__15226));
    CascadeMux I__2546 (
            .O(N__15235),
            .I(N__15223));
    CascadeMux I__2545 (
            .O(N__15232),
            .I(N__15220));
    CascadeMux I__2544 (
            .O(N__15229),
            .I(N__15217));
    CascadeMux I__2543 (
            .O(N__15226),
            .I(N__15214));
    InMux I__2542 (
            .O(N__15223),
            .I(N__15211));
    CascadeBuf I__2541 (
            .O(N__15220),
            .I(N__15208));
    CascadeBuf I__2540 (
            .O(N__15217),
            .I(N__15205));
    CascadeBuf I__2539 (
            .O(N__15214),
            .I(N__15202));
    LocalMux I__2538 (
            .O(N__15211),
            .I(N__15199));
    CascadeMux I__2537 (
            .O(N__15208),
            .I(N__15196));
    CascadeMux I__2536 (
            .O(N__15205),
            .I(N__15193));
    CascadeMux I__2535 (
            .O(N__15202),
            .I(N__15190));
    Span4Mux_s1_v I__2534 (
            .O(N__15199),
            .I(N__15186));
    InMux I__2533 (
            .O(N__15196),
            .I(N__15183));
    CascadeBuf I__2532 (
            .O(N__15193),
            .I(N__15180));
    InMux I__2531 (
            .O(N__15190),
            .I(N__15177));
    InMux I__2530 (
            .O(N__15189),
            .I(N__15174));
    Span4Mux_s2_h I__2529 (
            .O(N__15186),
            .I(N__15169));
    LocalMux I__2528 (
            .O(N__15183),
            .I(N__15169));
    CascadeMux I__2527 (
            .O(N__15180),
            .I(N__15166));
    LocalMux I__2526 (
            .O(N__15177),
            .I(N__15163));
    LocalMux I__2525 (
            .O(N__15174),
            .I(N__15158));
    Span4Mux_h I__2524 (
            .O(N__15169),
            .I(N__15158));
    InMux I__2523 (
            .O(N__15166),
            .I(N__15155));
    Span4Mux_s1_v I__2522 (
            .O(N__15163),
            .I(N__15148));
    Span4Mux_h I__2521 (
            .O(N__15158),
            .I(N__15148));
    LocalMux I__2520 (
            .O(N__15155),
            .I(N__15148));
    Span4Mux_v I__2519 (
            .O(N__15148),
            .I(N__15145));
    Span4Mux_v I__2518 (
            .O(N__15145),
            .I(N__15142));
    Odrv4 I__2517 (
            .O(N__15142),
            .I(addr_out_2));
    InMux I__2516 (
            .O(N__15139),
            .I(N__15136));
    LocalMux I__2515 (
            .O(N__15136),
            .I(N__15133));
    Odrv12 I__2514 (
            .O(N__15133),
            .I(\sb_translator_1.addr_out_RNO_0Z0Z_3 ));
    CascadeMux I__2513 (
            .O(N__15130),
            .I(N__15125));
    CascadeMux I__2512 (
            .O(N__15129),
            .I(N__15121));
    CascadeMux I__2511 (
            .O(N__15128),
            .I(N__15118));
    CascadeBuf I__2510 (
            .O(N__15125),
            .I(N__15115));
    CascadeMux I__2509 (
            .O(N__15124),
            .I(N__15112));
    CascadeBuf I__2508 (
            .O(N__15121),
            .I(N__15109));
    CascadeBuf I__2507 (
            .O(N__15118),
            .I(N__15106));
    CascadeMux I__2506 (
            .O(N__15115),
            .I(N__15103));
    CascadeBuf I__2505 (
            .O(N__15112),
            .I(N__15100));
    CascadeMux I__2504 (
            .O(N__15109),
            .I(N__15097));
    CascadeMux I__2503 (
            .O(N__15106),
            .I(N__15094));
    CascadeBuf I__2502 (
            .O(N__15103),
            .I(N__15091));
    CascadeMux I__2501 (
            .O(N__15100),
            .I(N__15088));
    CascadeBuf I__2500 (
            .O(N__15097),
            .I(N__15085));
    CascadeBuf I__2499 (
            .O(N__15094),
            .I(N__15082));
    CascadeMux I__2498 (
            .O(N__15091),
            .I(N__15079));
    CascadeBuf I__2497 (
            .O(N__15088),
            .I(N__15076));
    CascadeMux I__2496 (
            .O(N__15085),
            .I(N__15073));
    CascadeMux I__2495 (
            .O(N__15082),
            .I(N__15070));
    CascadeBuf I__2494 (
            .O(N__15079),
            .I(N__15067));
    CascadeMux I__2493 (
            .O(N__15076),
            .I(N__15064));
    CascadeBuf I__2492 (
            .O(N__15073),
            .I(N__15061));
    CascadeBuf I__2491 (
            .O(N__15070),
            .I(N__15058));
    CascadeMux I__2490 (
            .O(N__15067),
            .I(N__15055));
    CascadeBuf I__2489 (
            .O(N__15064),
            .I(N__15052));
    CascadeMux I__2488 (
            .O(N__15061),
            .I(N__15049));
    CascadeMux I__2487 (
            .O(N__15058),
            .I(N__15046));
    CascadeBuf I__2486 (
            .O(N__15055),
            .I(N__15043));
    CascadeMux I__2485 (
            .O(N__15052),
            .I(N__15040));
    CascadeBuf I__2484 (
            .O(N__15049),
            .I(N__15037));
    CascadeBuf I__2483 (
            .O(N__15046),
            .I(N__15034));
    CascadeMux I__2482 (
            .O(N__15043),
            .I(N__15031));
    CascadeBuf I__2481 (
            .O(N__15040),
            .I(N__15028));
    CascadeMux I__2480 (
            .O(N__15037),
            .I(N__15025));
    CascadeMux I__2479 (
            .O(N__15034),
            .I(N__15022));
    CascadeBuf I__2478 (
            .O(N__15031),
            .I(N__15019));
    CascadeMux I__2477 (
            .O(N__15028),
            .I(N__15016));
    CascadeBuf I__2476 (
            .O(N__15025),
            .I(N__15013));
    CascadeBuf I__2475 (
            .O(N__15022),
            .I(N__15010));
    CascadeMux I__2474 (
            .O(N__15019),
            .I(N__15007));
    CascadeBuf I__2473 (
            .O(N__15016),
            .I(N__15004));
    CascadeMux I__2472 (
            .O(N__15013),
            .I(N__15001));
    CascadeMux I__2471 (
            .O(N__15010),
            .I(N__14998));
    CascadeBuf I__2470 (
            .O(N__15007),
            .I(N__14995));
    CascadeMux I__2469 (
            .O(N__15004),
            .I(N__14992));
    CascadeBuf I__2468 (
            .O(N__15001),
            .I(N__14989));
    CascadeBuf I__2467 (
            .O(N__14998),
            .I(N__14986));
    CascadeMux I__2466 (
            .O(N__14995),
            .I(N__14983));
    CascadeBuf I__2465 (
            .O(N__14992),
            .I(N__14980));
    CascadeMux I__2464 (
            .O(N__14989),
            .I(N__14977));
    CascadeMux I__2463 (
            .O(N__14986),
            .I(N__14974));
    InMux I__2462 (
            .O(N__14983),
            .I(N__14970));
    CascadeMux I__2461 (
            .O(N__14980),
            .I(N__14967));
    InMux I__2460 (
            .O(N__14977),
            .I(N__14964));
    InMux I__2459 (
            .O(N__14974),
            .I(N__14961));
    InMux I__2458 (
            .O(N__14973),
            .I(N__14958));
    LocalMux I__2457 (
            .O(N__14970),
            .I(N__14955));
    InMux I__2456 (
            .O(N__14967),
            .I(N__14952));
    LocalMux I__2455 (
            .O(N__14964),
            .I(N__14949));
    LocalMux I__2454 (
            .O(N__14961),
            .I(N__14946));
    LocalMux I__2453 (
            .O(N__14958),
            .I(N__14941));
    Span4Mux_h I__2452 (
            .O(N__14955),
            .I(N__14941));
    LocalMux I__2451 (
            .O(N__14952),
            .I(N__14938));
    Span4Mux_h I__2450 (
            .O(N__14949),
            .I(N__14933));
    Span4Mux_h I__2449 (
            .O(N__14946),
            .I(N__14933));
    Span4Mux_h I__2448 (
            .O(N__14941),
            .I(N__14928));
    Span4Mux_h I__2447 (
            .O(N__14938),
            .I(N__14928));
    Span4Mux_v I__2446 (
            .O(N__14933),
            .I(N__14925));
    Span4Mux_v I__2445 (
            .O(N__14928),
            .I(N__14922));
    Span4Mux_v I__2444 (
            .O(N__14925),
            .I(N__14919));
    Span4Mux_v I__2443 (
            .O(N__14922),
            .I(N__14916));
    Odrv4 I__2442 (
            .O(N__14919),
            .I(addr_out_3));
    Odrv4 I__2441 (
            .O(N__14916),
            .I(addr_out_3));
    CascadeMux I__2440 (
            .O(N__14911),
            .I(N__14908));
    CascadeBuf I__2439 (
            .O(N__14908),
            .I(N__14902));
    CascadeMux I__2438 (
            .O(N__14907),
            .I(N__14899));
    CascadeMux I__2437 (
            .O(N__14906),
            .I(N__14896));
    CascadeMux I__2436 (
            .O(N__14905),
            .I(N__14893));
    CascadeMux I__2435 (
            .O(N__14902),
            .I(N__14890));
    CascadeBuf I__2434 (
            .O(N__14899),
            .I(N__14887));
    CascadeBuf I__2433 (
            .O(N__14896),
            .I(N__14884));
    CascadeBuf I__2432 (
            .O(N__14893),
            .I(N__14881));
    CascadeBuf I__2431 (
            .O(N__14890),
            .I(N__14878));
    CascadeMux I__2430 (
            .O(N__14887),
            .I(N__14875));
    CascadeMux I__2429 (
            .O(N__14884),
            .I(N__14872));
    CascadeMux I__2428 (
            .O(N__14881),
            .I(N__14869));
    CascadeMux I__2427 (
            .O(N__14878),
            .I(N__14866));
    CascadeBuf I__2426 (
            .O(N__14875),
            .I(N__14863));
    CascadeBuf I__2425 (
            .O(N__14872),
            .I(N__14860));
    CascadeBuf I__2424 (
            .O(N__14869),
            .I(N__14857));
    CascadeBuf I__2423 (
            .O(N__14866),
            .I(N__14854));
    CascadeMux I__2422 (
            .O(N__14863),
            .I(N__14851));
    CascadeMux I__2421 (
            .O(N__14860),
            .I(N__14848));
    CascadeMux I__2420 (
            .O(N__14857),
            .I(N__14845));
    CascadeMux I__2419 (
            .O(N__14854),
            .I(N__14842));
    CascadeBuf I__2418 (
            .O(N__14851),
            .I(N__14839));
    CascadeBuf I__2417 (
            .O(N__14848),
            .I(N__14836));
    CascadeBuf I__2416 (
            .O(N__14845),
            .I(N__14833));
    CascadeBuf I__2415 (
            .O(N__14842),
            .I(N__14830));
    CascadeMux I__2414 (
            .O(N__14839),
            .I(N__14827));
    CascadeMux I__2413 (
            .O(N__14836),
            .I(N__14824));
    CascadeMux I__2412 (
            .O(N__14833),
            .I(N__14821));
    CascadeMux I__2411 (
            .O(N__14830),
            .I(N__14818));
    CascadeBuf I__2410 (
            .O(N__14827),
            .I(N__14815));
    CascadeBuf I__2409 (
            .O(N__14824),
            .I(N__14812));
    CascadeBuf I__2408 (
            .O(N__14821),
            .I(N__14809));
    CascadeBuf I__2407 (
            .O(N__14818),
            .I(N__14806));
    CascadeMux I__2406 (
            .O(N__14815),
            .I(N__14803));
    CascadeMux I__2405 (
            .O(N__14812),
            .I(N__14800));
    CascadeMux I__2404 (
            .O(N__14809),
            .I(N__14797));
    CascadeMux I__2403 (
            .O(N__14806),
            .I(N__14794));
    CascadeBuf I__2402 (
            .O(N__14803),
            .I(N__14791));
    CascadeBuf I__2401 (
            .O(N__14800),
            .I(N__14788));
    CascadeBuf I__2400 (
            .O(N__14797),
            .I(N__14785));
    CascadeBuf I__2399 (
            .O(N__14794),
            .I(N__14782));
    CascadeMux I__2398 (
            .O(N__14791),
            .I(N__14779));
    CascadeMux I__2397 (
            .O(N__14788),
            .I(N__14776));
    CascadeMux I__2396 (
            .O(N__14785),
            .I(N__14773));
    CascadeMux I__2395 (
            .O(N__14782),
            .I(N__14770));
    CascadeBuf I__2394 (
            .O(N__14779),
            .I(N__14766));
    CascadeBuf I__2393 (
            .O(N__14776),
            .I(N__14763));
    CascadeBuf I__2392 (
            .O(N__14773),
            .I(N__14760));
    InMux I__2391 (
            .O(N__14770),
            .I(N__14757));
    InMux I__2390 (
            .O(N__14769),
            .I(N__14754));
    CascadeMux I__2389 (
            .O(N__14766),
            .I(N__14751));
    CascadeMux I__2388 (
            .O(N__14763),
            .I(N__14748));
    CascadeMux I__2387 (
            .O(N__14760),
            .I(N__14745));
    LocalMux I__2386 (
            .O(N__14757),
            .I(N__14742));
    LocalMux I__2385 (
            .O(N__14754),
            .I(N__14739));
    InMux I__2384 (
            .O(N__14751),
            .I(N__14736));
    InMux I__2383 (
            .O(N__14748),
            .I(N__14733));
    InMux I__2382 (
            .O(N__14745),
            .I(N__14730));
    Span4Mux_s1_v I__2381 (
            .O(N__14742),
            .I(N__14727));
    Span4Mux_h I__2380 (
            .O(N__14739),
            .I(N__14722));
    LocalMux I__2379 (
            .O(N__14736),
            .I(N__14722));
    LocalMux I__2378 (
            .O(N__14733),
            .I(N__14717));
    LocalMux I__2377 (
            .O(N__14730),
            .I(N__14717));
    Span4Mux_v I__2376 (
            .O(N__14727),
            .I(N__14712));
    Span4Mux_v I__2375 (
            .O(N__14722),
            .I(N__14712));
    Span12Mux_s9_v I__2374 (
            .O(N__14717),
            .I(N__14709));
    Span4Mux_v I__2373 (
            .O(N__14712),
            .I(N__14706));
    Odrv12 I__2372 (
            .O(N__14709),
            .I(addr_out_4));
    Odrv4 I__2371 (
            .O(N__14706),
            .I(addr_out_4));
    CascadeMux I__2370 (
            .O(N__14701),
            .I(\sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_ ));
    InMux I__2369 (
            .O(N__14698),
            .I(N__14695));
    LocalMux I__2368 (
            .O(N__14695),
            .I(miso_data_in_13));
    InMux I__2367 (
            .O(N__14692),
            .I(N__14689));
    LocalMux I__2366 (
            .O(N__14689),
            .I(miso_data_in_14));
    InMux I__2365 (
            .O(N__14686),
            .I(N__14683));
    LocalMux I__2364 (
            .O(N__14683),
            .I(miso_data_in_15));
    InMux I__2363 (
            .O(N__14680),
            .I(N__14677));
    LocalMux I__2362 (
            .O(N__14677),
            .I(miso_data_in_16));
    InMux I__2361 (
            .O(N__14674),
            .I(N__14671));
    LocalMux I__2360 (
            .O(N__14671),
            .I(N__14668));
    Span4Mux_h I__2359 (
            .O(N__14668),
            .I(N__14664));
    CascadeMux I__2358 (
            .O(N__14667),
            .I(N__14661));
    Span4Mux_h I__2357 (
            .O(N__14664),
            .I(N__14658));
    InMux I__2356 (
            .O(N__14661),
            .I(N__14655));
    Odrv4 I__2355 (
            .O(N__14658),
            .I(\sb_translator_1.instr_tmpZ0Z_17 ));
    LocalMux I__2354 (
            .O(N__14655),
            .I(\sb_translator_1.instr_tmpZ0Z_17 ));
    InMux I__2353 (
            .O(N__14650),
            .I(N__14647));
    LocalMux I__2352 (
            .O(N__14647),
            .I(miso_data_in_17));
    InMux I__2351 (
            .O(N__14644),
            .I(N__14640));
    InMux I__2350 (
            .O(N__14643),
            .I(N__14637));
    LocalMux I__2349 (
            .O(N__14640),
            .I(mosi_data_out_11));
    LocalMux I__2348 (
            .O(N__14637),
            .I(mosi_data_out_11));
    InMux I__2347 (
            .O(N__14632),
            .I(N__14629));
    LocalMux I__2346 (
            .O(N__14629),
            .I(N__14625));
    InMux I__2345 (
            .O(N__14628),
            .I(N__14621));
    Span4Mux_h I__2344 (
            .O(N__14625),
            .I(N__14618));
    InMux I__2343 (
            .O(N__14624),
            .I(N__14615));
    LocalMux I__2342 (
            .O(N__14621),
            .I(N__14612));
    Odrv4 I__2341 (
            .O(N__14618),
            .I(\sb_translator_1.cntZ0Z_3 ));
    LocalMux I__2340 (
            .O(N__14615),
            .I(\sb_translator_1.cntZ0Z_3 ));
    Odrv4 I__2339 (
            .O(N__14612),
            .I(\sb_translator_1.cntZ0Z_3 ));
    InMux I__2338 (
            .O(N__14605),
            .I(N__14601));
    InMux I__2337 (
            .O(N__14604),
            .I(N__14598));
    LocalMux I__2336 (
            .O(N__14601),
            .I(mosi_data_out_13));
    LocalMux I__2335 (
            .O(N__14598),
            .I(mosi_data_out_13));
    InMux I__2334 (
            .O(N__14593),
            .I(N__14590));
    LocalMux I__2333 (
            .O(N__14590),
            .I(N__14586));
    InMux I__2332 (
            .O(N__14589),
            .I(N__14582));
    Span4Mux_v I__2331 (
            .O(N__14586),
            .I(N__14579));
    InMux I__2330 (
            .O(N__14585),
            .I(N__14576));
    LocalMux I__2329 (
            .O(N__14582),
            .I(N__14573));
    Odrv4 I__2328 (
            .O(N__14579),
            .I(\sb_translator_1.cntZ0Z_5 ));
    LocalMux I__2327 (
            .O(N__14576),
            .I(\sb_translator_1.cntZ0Z_5 ));
    Odrv4 I__2326 (
            .O(N__14573),
            .I(\sb_translator_1.cntZ0Z_5 ));
    CascadeMux I__2325 (
            .O(N__14566),
            .I(N__14563));
    InMux I__2324 (
            .O(N__14563),
            .I(N__14560));
    LocalMux I__2323 (
            .O(N__14560),
            .I(N__14557));
    Span4Mux_h I__2322 (
            .O(N__14557),
            .I(N__14554));
    Odrv4 I__2321 (
            .O(N__14554),
            .I(\spi_slave_1.miso_data_outZ0Z_17 ));
    CEMux I__2320 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__2319 (
            .O(N__14548),
            .I(N__14543));
    CEMux I__2318 (
            .O(N__14547),
            .I(N__14540));
    CEMux I__2317 (
            .O(N__14546),
            .I(N__14536));
    Span4Mux_h I__2316 (
            .O(N__14543),
            .I(N__14531));
    LocalMux I__2315 (
            .O(N__14540),
            .I(N__14531));
    CEMux I__2314 (
            .O(N__14539),
            .I(N__14528));
    LocalMux I__2313 (
            .O(N__14536),
            .I(N__14525));
    Span4Mux_v I__2312 (
            .O(N__14531),
            .I(N__14520));
    LocalMux I__2311 (
            .O(N__14528),
            .I(N__14520));
    Span4Mux_v I__2310 (
            .O(N__14525),
            .I(N__14517));
    Span4Mux_h I__2309 (
            .O(N__14520),
            .I(N__14514));
    Odrv4 I__2308 (
            .O(N__14517),
            .I(\spi_slave_1.bitcnt_tx_0_sqmuxa ));
    Odrv4 I__2307 (
            .O(N__14514),
            .I(\spi_slave_1.bitcnt_tx_0_sqmuxa ));
    InMux I__2306 (
            .O(N__14509),
            .I(N__14506));
    LocalMux I__2305 (
            .O(N__14506),
            .I(miso_data_in_10));
    InMux I__2304 (
            .O(N__14503),
            .I(N__14500));
    LocalMux I__2303 (
            .O(N__14500),
            .I(miso_data_in_11));
    InMux I__2302 (
            .O(N__14497),
            .I(N__14494));
    LocalMux I__2301 (
            .O(N__14494),
            .I(miso_data_in_12));
    CascadeMux I__2300 (
            .O(N__14491),
            .I(\demux.N_236_cascade_ ));
    CascadeMux I__2299 (
            .O(N__14488),
            .I(\demux.N_235_cascade_ ));
    InMux I__2298 (
            .O(N__14485),
            .I(N__14479));
    InMux I__2297 (
            .O(N__14484),
            .I(N__14479));
    LocalMux I__2296 (
            .O(N__14479),
            .I(N__14473));
    InMux I__2295 (
            .O(N__14478),
            .I(N__14463));
    InMux I__2294 (
            .O(N__14477),
            .I(N__14463));
    InMux I__2293 (
            .O(N__14476),
            .I(N__14463));
    Span4Mux_h I__2292 (
            .O(N__14473),
            .I(N__14460));
    InMux I__2291 (
            .O(N__14472),
            .I(N__14453));
    InMux I__2290 (
            .O(N__14471),
            .I(N__14453));
    InMux I__2289 (
            .O(N__14470),
            .I(N__14453));
    LocalMux I__2288 (
            .O(N__14463),
            .I(N__14450));
    Odrv4 I__2287 (
            .O(N__14460),
            .I(\demux.N_424_i_0_a2Z0Z_6 ));
    LocalMux I__2286 (
            .O(N__14453),
            .I(\demux.N_424_i_0_a2Z0Z_6 ));
    Odrv12 I__2285 (
            .O(N__14450),
            .I(\demux.N_424_i_0_a2Z0Z_6 ));
    CascadeMux I__2284 (
            .O(N__14443),
            .I(N__14439));
    InMux I__2283 (
            .O(N__14442),
            .I(N__14425));
    InMux I__2282 (
            .O(N__14439),
            .I(N__14425));
    InMux I__2281 (
            .O(N__14438),
            .I(N__14425));
    InMux I__2280 (
            .O(N__14437),
            .I(N__14425));
    InMux I__2279 (
            .O(N__14436),
            .I(N__14425));
    LocalMux I__2278 (
            .O(N__14425),
            .I(N__14422));
    Odrv4 I__2277 (
            .O(N__14422),
            .I(ram_sel_6));
    InMux I__2276 (
            .O(N__14419),
            .I(N__14404));
    InMux I__2275 (
            .O(N__14418),
            .I(N__14404));
    InMux I__2274 (
            .O(N__14417),
            .I(N__14404));
    InMux I__2273 (
            .O(N__14416),
            .I(N__14404));
    InMux I__2272 (
            .O(N__14415),
            .I(N__14404));
    LocalMux I__2271 (
            .O(N__14404),
            .I(N__14401));
    Odrv4 I__2270 (
            .O(N__14401),
            .I(ram_sel_9));
    InMux I__2269 (
            .O(N__14398),
            .I(N__14395));
    LocalMux I__2268 (
            .O(N__14395),
            .I(N__14392));
    Span4Mux_s3_v I__2267 (
            .O(N__14392),
            .I(N__14389));
    Span4Mux_h I__2266 (
            .O(N__14389),
            .I(N__14386));
    Odrv4 I__2265 (
            .O(N__14386),
            .I(miso_data_in_9));
    InMux I__2264 (
            .O(N__14383),
            .I(N__14380));
    LocalMux I__2263 (
            .O(N__14380),
            .I(N__14377));
    Span4Mux_h I__2262 (
            .O(N__14377),
            .I(N__14374));
    Odrv4 I__2261 (
            .O(N__14374),
            .I(demux_data_in_56));
    InMux I__2260 (
            .O(N__14371),
            .I(N__14368));
    LocalMux I__2259 (
            .O(N__14368),
            .I(\demux.N_424_i_0_a3Z0Z_1 ));
    InMux I__2258 (
            .O(N__14365),
            .I(N__14356));
    InMux I__2257 (
            .O(N__14364),
            .I(N__14356));
    InMux I__2256 (
            .O(N__14363),
            .I(N__14356));
    LocalMux I__2255 (
            .O(N__14356),
            .I(N__14353));
    Odrv4 I__2254 (
            .O(N__14353),
            .I(\sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9 ));
    CascadeMux I__2253 (
            .O(N__14350),
            .I(N__14347));
    InMux I__2252 (
            .O(N__14347),
            .I(N__14338));
    InMux I__2251 (
            .O(N__14346),
            .I(N__14333));
    InMux I__2250 (
            .O(N__14345),
            .I(N__14333));
    InMux I__2249 (
            .O(N__14344),
            .I(N__14324));
    InMux I__2248 (
            .O(N__14343),
            .I(N__14324));
    InMux I__2247 (
            .O(N__14342),
            .I(N__14324));
    InMux I__2246 (
            .O(N__14341),
            .I(N__14324));
    LocalMux I__2245 (
            .O(N__14338),
            .I(N__14319));
    LocalMux I__2244 (
            .O(N__14333),
            .I(N__14319));
    LocalMux I__2243 (
            .O(N__14324),
            .I(\sb_translator_1.state_RNIHS98Z0Z_0 ));
    Odrv4 I__2242 (
            .O(N__14319),
            .I(\sb_translator_1.state_RNIHS98Z0Z_0 ));
    InMux I__2241 (
            .O(N__14314),
            .I(N__14299));
    InMux I__2240 (
            .O(N__14313),
            .I(N__14299));
    InMux I__2239 (
            .O(N__14312),
            .I(N__14299));
    InMux I__2238 (
            .O(N__14311),
            .I(N__14299));
    InMux I__2237 (
            .O(N__14310),
            .I(N__14299));
    LocalMux I__2236 (
            .O(N__14299),
            .I(N__14296));
    Span4Mux_v I__2235 (
            .O(N__14296),
            .I(N__14292));
    InMux I__2234 (
            .O(N__14295),
            .I(N__14289));
    Odrv4 I__2233 (
            .O(N__14292),
            .I(\sb_translator_1.state_RNIHS98_0Z0Z_0 ));
    LocalMux I__2232 (
            .O(N__14289),
            .I(\sb_translator_1.state_RNIHS98_0Z0Z_0 ));
    CascadeMux I__2231 (
            .O(N__14284),
            .I(N__14278));
    InMux I__2230 (
            .O(N__14283),
            .I(N__14275));
    InMux I__2229 (
            .O(N__14282),
            .I(N__14272));
    CascadeMux I__2228 (
            .O(N__14281),
            .I(N__14269));
    InMux I__2227 (
            .O(N__14278),
            .I(N__14266));
    LocalMux I__2226 (
            .O(N__14275),
            .I(N__14261));
    LocalMux I__2225 (
            .O(N__14272),
            .I(N__14261));
    InMux I__2224 (
            .O(N__14269),
            .I(N__14258));
    LocalMux I__2223 (
            .O(N__14266),
            .I(N__14255));
    Span4Mux_h I__2222 (
            .O(N__14261),
            .I(N__14252));
    LocalMux I__2221 (
            .O(N__14258),
            .I(N__14249));
    Span4Mux_h I__2220 (
            .O(N__14255),
            .I(N__14246));
    Span4Mux_s2_h I__2219 (
            .O(N__14252),
            .I(N__14243));
    Span4Mux_h I__2218 (
            .O(N__14249),
            .I(N__14240));
    Odrv4 I__2217 (
            .O(N__14246),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9 ));
    Odrv4 I__2216 (
            .O(N__14243),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9 ));
    Odrv4 I__2215 (
            .O(N__14240),
            .I(\sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9 ));
    CascadeMux I__2214 (
            .O(N__14233),
            .I(N__14229));
    InMux I__2213 (
            .O(N__14232),
            .I(N__14224));
    InMux I__2212 (
            .O(N__14229),
            .I(N__14224));
    LocalMux I__2211 (
            .O(N__14224),
            .I(N__14221));
    Odrv4 I__2210 (
            .O(N__14221),
            .I(\sb_translator_1.N_1089 ));
    CascadeMux I__2209 (
            .O(N__14218),
            .I(\sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_ ));
    InMux I__2208 (
            .O(N__14215),
            .I(N__14212));
    LocalMux I__2207 (
            .O(N__14212),
            .I(N__14209));
    Span4Mux_h I__2206 (
            .O(N__14209),
            .I(N__14206));
    Span4Mux_v I__2205 (
            .O(N__14206),
            .I(N__14203));
    Odrv4 I__2204 (
            .O(N__14203),
            .I(demux_data_in_74));
    CascadeMux I__2203 (
            .O(N__14200),
            .I(N__14197));
    InMux I__2202 (
            .O(N__14197),
            .I(N__14194));
    LocalMux I__2201 (
            .O(N__14194),
            .I(N__14191));
    Span4Mux_v I__2200 (
            .O(N__14191),
            .I(N__14188));
    Span4Mux_h I__2199 (
            .O(N__14188),
            .I(N__14185));
    Odrv4 I__2198 (
            .O(N__14185),
            .I(demux_data_in_82));
    InMux I__2197 (
            .O(N__14182),
            .I(N__14179));
    LocalMux I__2196 (
            .O(N__14179),
            .I(N__14176));
    Span4Mux_h I__2195 (
            .O(N__14176),
            .I(N__14173));
    Odrv4 I__2194 (
            .O(N__14173),
            .I(demux_data_in_50));
    CascadeMux I__2193 (
            .O(N__14170),
            .I(\demux.N_422_i_0_o2Z0Z_6_cascade_ ));
    InMux I__2192 (
            .O(N__14167),
            .I(N__14164));
    LocalMux I__2191 (
            .O(N__14164),
            .I(N__14161));
    Span4Mux_h I__2190 (
            .O(N__14161),
            .I(N__14158));
    Span4Mux_v I__2189 (
            .O(N__14158),
            .I(N__14155));
    Odrv4 I__2188 (
            .O(N__14155),
            .I(demux_data_in_73));
    CascadeMux I__2187 (
            .O(N__14152),
            .I(N__14149));
    InMux I__2186 (
            .O(N__14149),
            .I(N__14146));
    LocalMux I__2185 (
            .O(N__14146),
            .I(N__14143));
    Span12Mux_s10_h I__2184 (
            .O(N__14143),
            .I(N__14140));
    Odrv12 I__2183 (
            .O(N__14140),
            .I(demux_data_in_81));
    InMux I__2182 (
            .O(N__14137),
            .I(N__14134));
    LocalMux I__2181 (
            .O(N__14134),
            .I(N__14131));
    Span4Mux_v I__2180 (
            .O(N__14131),
            .I(N__14128));
    Odrv4 I__2179 (
            .O(N__14128),
            .I(demux_data_in_49));
    CascadeMux I__2178 (
            .O(N__14125),
            .I(\demux.N_423_i_0_o2Z0Z_6_cascade_ ));
    InMux I__2177 (
            .O(N__14122),
            .I(N__14119));
    LocalMux I__2176 (
            .O(N__14119),
            .I(\demux.N_423_i_0_a3Z0Z_1 ));
    InMux I__2175 (
            .O(N__14116),
            .I(N__14113));
    LocalMux I__2174 (
            .O(N__14113),
            .I(N__14110));
    Span4Mux_h I__2173 (
            .O(N__14110),
            .I(N__14107));
    Odrv4 I__2172 (
            .O(N__14107),
            .I(demux_data_in_58));
    InMux I__2171 (
            .O(N__14104),
            .I(N__14101));
    LocalMux I__2170 (
            .O(N__14101),
            .I(\demux.N_422_i_0_a3Z0Z_1 ));
    InMux I__2169 (
            .O(N__14098),
            .I(N__14095));
    LocalMux I__2168 (
            .O(N__14095),
            .I(N__14092));
    Span4Mux_v I__2167 (
            .O(N__14092),
            .I(N__14089));
    Span4Mux_h I__2166 (
            .O(N__14089),
            .I(N__14086));
    Odrv4 I__2165 (
            .O(N__14086),
            .I(demux_data_in_80));
    InMux I__2164 (
            .O(N__14083),
            .I(N__14080));
    LocalMux I__2163 (
            .O(N__14080),
            .I(N__14077));
    Span12Mux_s10_h I__2162 (
            .O(N__14077),
            .I(N__14074));
    Odrv12 I__2161 (
            .O(N__14074),
            .I(demux_data_in_72));
    InMux I__2160 (
            .O(N__14071),
            .I(N__14068));
    LocalMux I__2159 (
            .O(N__14068),
            .I(N__14065));
    Span4Mux_h I__2158 (
            .O(N__14065),
            .I(N__14062));
    Span4Mux_s3_h I__2157 (
            .O(N__14062),
            .I(N__14059));
    Odrv4 I__2156 (
            .O(N__14059),
            .I(demux_data_in_48));
    CascadeMux I__2155 (
            .O(N__14056),
            .I(\demux.N_424_i_0_o2_6_cascade_ ));
    CascadeMux I__2154 (
            .O(N__14053),
            .I(N__14050));
    InMux I__2153 (
            .O(N__14050),
            .I(N__14043));
    InMux I__2152 (
            .O(N__14049),
            .I(N__14043));
    InMux I__2151 (
            .O(N__14048),
            .I(N__14040));
    LocalMux I__2150 (
            .O(N__14043),
            .I(\sb_translator_1.cnt_RNILAHE_0Z0Z_10 ));
    LocalMux I__2149 (
            .O(N__14040),
            .I(\sb_translator_1.cnt_RNILAHE_0Z0Z_10 ));
    CEMux I__2148 (
            .O(N__14035),
            .I(N__14032));
    LocalMux I__2147 (
            .O(N__14032),
            .I(N__14029));
    Span4Mux_h I__2146 (
            .O(N__14029),
            .I(N__14026));
    Span4Mux_h I__2145 (
            .O(N__14026),
            .I(N__14023));
    Sp12to4 I__2144 (
            .O(N__14023),
            .I(N__14020));
    Span12Mux_s6_v I__2143 (
            .O(N__14020),
            .I(N__14017));
    Odrv12 I__2142 (
            .O(N__14017),
            .I(ram_we_4));
    InMux I__2141 (
            .O(N__14014),
            .I(N__14002));
    InMux I__2140 (
            .O(N__14013),
            .I(N__14002));
    InMux I__2139 (
            .O(N__14012),
            .I(N__14002));
    InMux I__2138 (
            .O(N__14011),
            .I(N__14002));
    LocalMux I__2137 (
            .O(N__14002),
            .I(N__13999));
    Span4Mux_h I__2136 (
            .O(N__13999),
            .I(N__13996));
    Odrv4 I__2135 (
            .O(N__13996),
            .I(\sb_translator_1.cnt_RNIJ7EF_2Z0Z_9 ));
    InMux I__2134 (
            .O(N__13993),
            .I(N__13972));
    InMux I__2133 (
            .O(N__13992),
            .I(N__13972));
    InMux I__2132 (
            .O(N__13991),
            .I(N__13972));
    InMux I__2131 (
            .O(N__13990),
            .I(N__13972));
    InMux I__2130 (
            .O(N__13989),
            .I(N__13972));
    InMux I__2129 (
            .O(N__13988),
            .I(N__13972));
    InMux I__2128 (
            .O(N__13987),
            .I(N__13972));
    LocalMux I__2127 (
            .O(N__13972),
            .I(\sb_translator_1.state_RNI9ILJ_0Z0Z_0 ));
    CEMux I__2126 (
            .O(N__13969),
            .I(N__13966));
    LocalMux I__2125 (
            .O(N__13966),
            .I(N__13963));
    Span4Mux_v I__2124 (
            .O(N__13963),
            .I(N__13960));
    Sp12to4 I__2123 (
            .O(N__13960),
            .I(N__13957));
    Span12Mux_s7_v I__2122 (
            .O(N__13957),
            .I(N__13954));
    Odrv12 I__2121 (
            .O(N__13954),
            .I(ram_we_6));
    InMux I__2120 (
            .O(N__13951),
            .I(N__13948));
    LocalMux I__2119 (
            .O(N__13948),
            .I(N__13942));
    InMux I__2118 (
            .O(N__13947),
            .I(N__13935));
    InMux I__2117 (
            .O(N__13946),
            .I(N__13935));
    InMux I__2116 (
            .O(N__13945),
            .I(N__13935));
    Span4Mux_h I__2115 (
            .O(N__13942),
            .I(N__13932));
    LocalMux I__2114 (
            .O(N__13935),
            .I(N__13929));
    Odrv4 I__2113 (
            .O(N__13932),
            .I(\sb_translator_1.cnt_RNIJ7EF_1Z0Z_9 ));
    Odrv12 I__2112 (
            .O(N__13929),
            .I(\sb_translator_1.cnt_RNIJ7EF_1Z0Z_9 ));
    InMux I__2111 (
            .O(N__13924),
            .I(N__13915));
    InMux I__2110 (
            .O(N__13923),
            .I(N__13902));
    InMux I__2109 (
            .O(N__13922),
            .I(N__13902));
    InMux I__2108 (
            .O(N__13921),
            .I(N__13902));
    InMux I__2107 (
            .O(N__13920),
            .I(N__13902));
    InMux I__2106 (
            .O(N__13919),
            .I(N__13902));
    InMux I__2105 (
            .O(N__13918),
            .I(N__13902));
    LocalMux I__2104 (
            .O(N__13915),
            .I(\sb_translator_1.state_RNI9ILJZ0Z_0 ));
    LocalMux I__2103 (
            .O(N__13902),
            .I(\sb_translator_1.state_RNI9ILJZ0Z_0 ));
    CEMux I__2102 (
            .O(N__13897),
            .I(N__13894));
    LocalMux I__2101 (
            .O(N__13894),
            .I(N__13891));
    Span4Mux_s3_h I__2100 (
            .O(N__13891),
            .I(N__13888));
    Span4Mux_h I__2099 (
            .O(N__13888),
            .I(N__13885));
    Span4Mux_v I__2098 (
            .O(N__13885),
            .I(N__13882));
    Odrv4 I__2097 (
            .O(N__13882),
            .I(ram_we_1));
    CascadeMux I__2096 (
            .O(N__13879),
            .I(\sb_translator_1.N_1091_cascade_ ));
    CascadeMux I__2095 (
            .O(N__13876),
            .I(\sb_translator_1.N_1089_cascade_ ));
    CascadeMux I__2094 (
            .O(N__13873),
            .I(N__13869));
    InMux I__2093 (
            .O(N__13872),
            .I(N__13864));
    InMux I__2092 (
            .O(N__13869),
            .I(N__13864));
    LocalMux I__2091 (
            .O(N__13864),
            .I(\sb_translator_1.N_1091 ));
    InMux I__2090 (
            .O(N__13861),
            .I(N__13858));
    LocalMux I__2089 (
            .O(N__13858),
            .I(\sb_translator_1.instr_tmpZ1Z_5 ));
    InMux I__2088 (
            .O(N__13855),
            .I(N__13852));
    LocalMux I__2087 (
            .O(N__13852),
            .I(N__13849));
    Span4Mux_s1_v I__2086 (
            .O(N__13849),
            .I(N__13844));
    InMux I__2085 (
            .O(N__13848),
            .I(N__13841));
    InMux I__2084 (
            .O(N__13847),
            .I(N__13838));
    Odrv4 I__2083 (
            .O(N__13844),
            .I(mosi_data_out_5));
    LocalMux I__2082 (
            .O(N__13841),
            .I(mosi_data_out_5));
    LocalMux I__2081 (
            .O(N__13838),
            .I(mosi_data_out_5));
    InMux I__2080 (
            .O(N__13831),
            .I(N__13827));
    InMux I__2079 (
            .O(N__13830),
            .I(N__13819));
    LocalMux I__2078 (
            .O(N__13827),
            .I(N__13815));
    InMux I__2077 (
            .O(N__13826),
            .I(N__13812));
    InMux I__2076 (
            .O(N__13825),
            .I(N__13809));
    InMux I__2075 (
            .O(N__13824),
            .I(N__13806));
    InMux I__2074 (
            .O(N__13823),
            .I(N__13803));
    InMux I__2073 (
            .O(N__13822),
            .I(N__13799));
    LocalMux I__2072 (
            .O(N__13819),
            .I(N__13795));
    InMux I__2071 (
            .O(N__13818),
            .I(N__13792));
    Span4Mux_s3_v I__2070 (
            .O(N__13815),
            .I(N__13781));
    LocalMux I__2069 (
            .O(N__13812),
            .I(N__13781));
    LocalMux I__2068 (
            .O(N__13809),
            .I(N__13781));
    LocalMux I__2067 (
            .O(N__13806),
            .I(N__13776));
    LocalMux I__2066 (
            .O(N__13803),
            .I(N__13776));
    InMux I__2065 (
            .O(N__13802),
            .I(N__13773));
    LocalMux I__2064 (
            .O(N__13799),
            .I(N__13770));
    InMux I__2063 (
            .O(N__13798),
            .I(N__13767));
    Span4Mux_s3_h I__2062 (
            .O(N__13795),
            .I(N__13762));
    LocalMux I__2061 (
            .O(N__13792),
            .I(N__13762));
    InMux I__2060 (
            .O(N__13791),
            .I(N__13759));
    InMux I__2059 (
            .O(N__13790),
            .I(N__13756));
    InMux I__2058 (
            .O(N__13789),
            .I(N__13753));
    InMux I__2057 (
            .O(N__13788),
            .I(N__13750));
    Span4Mux_v I__2056 (
            .O(N__13781),
            .I(N__13743));
    Span4Mux_s2_v I__2055 (
            .O(N__13776),
            .I(N__13743));
    LocalMux I__2054 (
            .O(N__13773),
            .I(N__13743));
    Span4Mux_s0_v I__2053 (
            .O(N__13770),
            .I(N__13738));
    LocalMux I__2052 (
            .O(N__13767),
            .I(N__13738));
    Span4Mux_v I__2051 (
            .O(N__13762),
            .I(N__13731));
    LocalMux I__2050 (
            .O(N__13759),
            .I(N__13731));
    LocalMux I__2049 (
            .O(N__13756),
            .I(N__13731));
    LocalMux I__2048 (
            .O(N__13753),
            .I(N__13728));
    LocalMux I__2047 (
            .O(N__13750),
            .I(N__13725));
    Sp12to4 I__2046 (
            .O(N__13743),
            .I(N__13722));
    Span4Mux_v I__2045 (
            .O(N__13738),
            .I(N__13713));
    Span4Mux_v I__2044 (
            .O(N__13731),
            .I(N__13713));
    Span4Mux_s3_h I__2043 (
            .O(N__13728),
            .I(N__13713));
    Span4Mux_h I__2042 (
            .O(N__13725),
            .I(N__13713));
    Span12Mux_s5_v I__2041 (
            .O(N__13722),
            .I(N__13710));
    Span4Mux_h I__2040 (
            .O(N__13713),
            .I(N__13707));
    Odrv12 I__2039 (
            .O(N__13710),
            .I(ram_data_in_5));
    Odrv4 I__2038 (
            .O(N__13707),
            .I(ram_data_in_5));
    InMux I__2037 (
            .O(N__13702),
            .I(N__13699));
    LocalMux I__2036 (
            .O(N__13699),
            .I(N__13696));
    Odrv4 I__2035 (
            .O(N__13696),
            .I(\sb_translator_1.instr_tmpZ0Z_6 ));
    InMux I__2034 (
            .O(N__13693),
            .I(N__13690));
    LocalMux I__2033 (
            .O(N__13690),
            .I(N__13685));
    InMux I__2032 (
            .O(N__13689),
            .I(N__13682));
    InMux I__2031 (
            .O(N__13688),
            .I(N__13679));
    Odrv4 I__2030 (
            .O(N__13685),
            .I(mosi_data_out_6));
    LocalMux I__2029 (
            .O(N__13682),
            .I(mosi_data_out_6));
    LocalMux I__2028 (
            .O(N__13679),
            .I(mosi_data_out_6));
    InMux I__2027 (
            .O(N__13672),
            .I(N__13666));
    InMux I__2026 (
            .O(N__13671),
            .I(N__13659));
    InMux I__2025 (
            .O(N__13670),
            .I(N__13656));
    InMux I__2024 (
            .O(N__13669),
            .I(N__13652));
    LocalMux I__2023 (
            .O(N__13666),
            .I(N__13649));
    InMux I__2022 (
            .O(N__13665),
            .I(N__13646));
    InMux I__2021 (
            .O(N__13664),
            .I(N__13642));
    InMux I__2020 (
            .O(N__13663),
            .I(N__13639));
    InMux I__2019 (
            .O(N__13662),
            .I(N__13635));
    LocalMux I__2018 (
            .O(N__13659),
            .I(N__13631));
    LocalMux I__2017 (
            .O(N__13656),
            .I(N__13628));
    InMux I__2016 (
            .O(N__13655),
            .I(N__13625));
    LocalMux I__2015 (
            .O(N__13652),
            .I(N__13621));
    Span4Mux_h I__2014 (
            .O(N__13649),
            .I(N__13618));
    LocalMux I__2013 (
            .O(N__13646),
            .I(N__13615));
    InMux I__2012 (
            .O(N__13645),
            .I(N__13612));
    LocalMux I__2011 (
            .O(N__13642),
            .I(N__13606));
    LocalMux I__2010 (
            .O(N__13639),
            .I(N__13606));
    InMux I__2009 (
            .O(N__13638),
            .I(N__13603));
    LocalMux I__2008 (
            .O(N__13635),
            .I(N__13600));
    InMux I__2007 (
            .O(N__13634),
            .I(N__13597));
    Span4Mux_h I__2006 (
            .O(N__13631),
            .I(N__13594));
    Span4Mux_h I__2005 (
            .O(N__13628),
            .I(N__13591));
    LocalMux I__2004 (
            .O(N__13625),
            .I(N__13588));
    InMux I__2003 (
            .O(N__13624),
            .I(N__13585));
    Span4Mux_h I__2002 (
            .O(N__13621),
            .I(N__13582));
    Span4Mux_v I__2001 (
            .O(N__13618),
            .I(N__13577));
    Span4Mux_h I__2000 (
            .O(N__13615),
            .I(N__13577));
    LocalMux I__1999 (
            .O(N__13612),
            .I(N__13574));
    InMux I__1998 (
            .O(N__13611),
            .I(N__13571));
    Span4Mux_v I__1997 (
            .O(N__13606),
            .I(N__13566));
    LocalMux I__1996 (
            .O(N__13603),
            .I(N__13566));
    Span4Mux_s1_v I__1995 (
            .O(N__13600),
            .I(N__13561));
    LocalMux I__1994 (
            .O(N__13597),
            .I(N__13561));
    Span4Mux_v I__1993 (
            .O(N__13594),
            .I(N__13554));
    Span4Mux_v I__1992 (
            .O(N__13591),
            .I(N__13554));
    Span4Mux_h I__1991 (
            .O(N__13588),
            .I(N__13554));
    LocalMux I__1990 (
            .O(N__13585),
            .I(N__13551));
    Span4Mux_v I__1989 (
            .O(N__13582),
            .I(N__13544));
    Span4Mux_v I__1988 (
            .O(N__13577),
            .I(N__13544));
    Span4Mux_h I__1987 (
            .O(N__13574),
            .I(N__13544));
    LocalMux I__1986 (
            .O(N__13571),
            .I(N__13541));
    Span4Mux_v I__1985 (
            .O(N__13566),
            .I(N__13536));
    Span4Mux_v I__1984 (
            .O(N__13561),
            .I(N__13536));
    Span4Mux_h I__1983 (
            .O(N__13554),
            .I(N__13531));
    Span4Mux_h I__1982 (
            .O(N__13551),
            .I(N__13531));
    Span4Mux_h I__1981 (
            .O(N__13544),
            .I(N__13526));
    Span4Mux_h I__1980 (
            .O(N__13541),
            .I(N__13526));
    Odrv4 I__1979 (
            .O(N__13536),
            .I(ram_data_in_6));
    Odrv4 I__1978 (
            .O(N__13531),
            .I(ram_data_in_6));
    Odrv4 I__1977 (
            .O(N__13526),
            .I(ram_data_in_6));
    InMux I__1976 (
            .O(N__13519),
            .I(N__13516));
    LocalMux I__1975 (
            .O(N__13516),
            .I(\sb_translator_1.instr_tmpZ0Z_7 ));
    InMux I__1974 (
            .O(N__13513),
            .I(N__13510));
    LocalMux I__1973 (
            .O(N__13510),
            .I(N__13505));
    InMux I__1972 (
            .O(N__13509),
            .I(N__13502));
    InMux I__1971 (
            .O(N__13508),
            .I(N__13499));
    Odrv4 I__1970 (
            .O(N__13505),
            .I(mosi_data_out_7));
    LocalMux I__1969 (
            .O(N__13502),
            .I(mosi_data_out_7));
    LocalMux I__1968 (
            .O(N__13499),
            .I(mosi_data_out_7));
    InMux I__1967 (
            .O(N__13492),
            .I(N__13488));
    InMux I__1966 (
            .O(N__13491),
            .I(N__13481));
    LocalMux I__1965 (
            .O(N__13488),
            .I(N__13478));
    InMux I__1964 (
            .O(N__13487),
            .I(N__13473));
    InMux I__1963 (
            .O(N__13486),
            .I(N__13468));
    InMux I__1962 (
            .O(N__13485),
            .I(N__13465));
    InMux I__1961 (
            .O(N__13484),
            .I(N__13461));
    LocalMux I__1960 (
            .O(N__13481),
            .I(N__13457));
    Span4Mux_h I__1959 (
            .O(N__13478),
            .I(N__13454));
    InMux I__1958 (
            .O(N__13477),
            .I(N__13451));
    InMux I__1957 (
            .O(N__13476),
            .I(N__13447));
    LocalMux I__1956 (
            .O(N__13473),
            .I(N__13444));
    InMux I__1955 (
            .O(N__13472),
            .I(N__13441));
    InMux I__1954 (
            .O(N__13471),
            .I(N__13437));
    LocalMux I__1953 (
            .O(N__13468),
            .I(N__13432));
    LocalMux I__1952 (
            .O(N__13465),
            .I(N__13432));
    InMux I__1951 (
            .O(N__13464),
            .I(N__13429));
    LocalMux I__1950 (
            .O(N__13461),
            .I(N__13426));
    InMux I__1949 (
            .O(N__13460),
            .I(N__13423));
    Span4Mux_h I__1948 (
            .O(N__13457),
            .I(N__13420));
    Span4Mux_v I__1947 (
            .O(N__13454),
            .I(N__13415));
    LocalMux I__1946 (
            .O(N__13451),
            .I(N__13415));
    InMux I__1945 (
            .O(N__13450),
            .I(N__13412));
    LocalMux I__1944 (
            .O(N__13447),
            .I(N__13409));
    Span4Mux_h I__1943 (
            .O(N__13444),
            .I(N__13406));
    LocalMux I__1942 (
            .O(N__13441),
            .I(N__13403));
    InMux I__1941 (
            .O(N__13440),
            .I(N__13400));
    LocalMux I__1940 (
            .O(N__13437),
            .I(N__13397));
    Span4Mux_v I__1939 (
            .O(N__13432),
            .I(N__13392));
    LocalMux I__1938 (
            .O(N__13429),
            .I(N__13392));
    Span4Mux_s1_v I__1937 (
            .O(N__13426),
            .I(N__13387));
    LocalMux I__1936 (
            .O(N__13423),
            .I(N__13387));
    Span4Mux_v I__1935 (
            .O(N__13420),
            .I(N__13382));
    Span4Mux_h I__1934 (
            .O(N__13415),
            .I(N__13382));
    LocalMux I__1933 (
            .O(N__13412),
            .I(N__13379));
    Span4Mux_h I__1932 (
            .O(N__13409),
            .I(N__13376));
    Span4Mux_v I__1931 (
            .O(N__13406),
            .I(N__13371));
    Span4Mux_h I__1930 (
            .O(N__13403),
            .I(N__13371));
    LocalMux I__1929 (
            .O(N__13400),
            .I(N__13368));
    Span12Mux_s8_h I__1928 (
            .O(N__13397),
            .I(N__13365));
    Span4Mux_v I__1927 (
            .O(N__13392),
            .I(N__13360));
    Span4Mux_v I__1926 (
            .O(N__13387),
            .I(N__13360));
    Span4Mux_h I__1925 (
            .O(N__13382),
            .I(N__13355));
    Span4Mux_h I__1924 (
            .O(N__13379),
            .I(N__13355));
    Span4Mux_h I__1923 (
            .O(N__13376),
            .I(N__13348));
    Span4Mux_h I__1922 (
            .O(N__13371),
            .I(N__13348));
    Span4Mux_h I__1921 (
            .O(N__13368),
            .I(N__13348));
    Odrv12 I__1920 (
            .O(N__13365),
            .I(ram_data_in_7));
    Odrv4 I__1919 (
            .O(N__13360),
            .I(ram_data_in_7));
    Odrv4 I__1918 (
            .O(N__13355),
            .I(ram_data_in_7));
    Odrv4 I__1917 (
            .O(N__13348),
            .I(ram_data_in_7));
    CEMux I__1916 (
            .O(N__13339),
            .I(N__13336));
    LocalMux I__1915 (
            .O(N__13336),
            .I(N__13333));
    Span4Mux_s2_v I__1914 (
            .O(N__13333),
            .I(N__13330));
    Span4Mux_h I__1913 (
            .O(N__13330),
            .I(N__13327));
    Odrv4 I__1912 (
            .O(N__13327),
            .I(ram_we_0));
    CEMux I__1911 (
            .O(N__13324),
            .I(N__13321));
    LocalMux I__1910 (
            .O(N__13321),
            .I(N__13318));
    Span4Mux_s1_v I__1909 (
            .O(N__13318),
            .I(N__13315));
    Span4Mux_h I__1908 (
            .O(N__13315),
            .I(N__13312));
    Span4Mux_v I__1907 (
            .O(N__13312),
            .I(N__13309));
    Odrv4 I__1906 (
            .O(N__13309),
            .I(ram_we_2));
    CascadeMux I__1905 (
            .O(N__13306),
            .I(N__13303));
    InMux I__1904 (
            .O(N__13303),
            .I(N__13296));
    InMux I__1903 (
            .O(N__13302),
            .I(N__13296));
    InMux I__1902 (
            .O(N__13301),
            .I(N__13293));
    LocalMux I__1901 (
            .O(N__13296),
            .I(\sb_translator_1.cnt_RNILAHE_1Z0Z_10 ));
    LocalMux I__1900 (
            .O(N__13293),
            .I(\sb_translator_1.cnt_RNILAHE_1Z0Z_10 ));
    CEMux I__1899 (
            .O(N__13288),
            .I(N__13285));
    LocalMux I__1898 (
            .O(N__13285),
            .I(N__13282));
    Span4Mux_s3_v I__1897 (
            .O(N__13282),
            .I(N__13279));
    Span4Mux_s3_h I__1896 (
            .O(N__13279),
            .I(N__13276));
    Span4Mux_h I__1895 (
            .O(N__13276),
            .I(N__13273));
    Odrv4 I__1894 (
            .O(N__13273),
            .I(ram_we_10));
    CEMux I__1893 (
            .O(N__13270),
            .I(N__13267));
    LocalMux I__1892 (
            .O(N__13267),
            .I(N__13264));
    Span4Mux_h I__1891 (
            .O(N__13264),
            .I(N__13261));
    Span4Mux_v I__1890 (
            .O(N__13261),
            .I(N__13258));
    Odrv4 I__1889 (
            .O(N__13258),
            .I(ram_we_8));
    CascadeMux I__1888 (
            .O(N__13255),
            .I(N__13251));
    InMux I__1887 (
            .O(N__13254),
            .I(N__13243));
    InMux I__1886 (
            .O(N__13251),
            .I(N__13243));
    InMux I__1885 (
            .O(N__13250),
            .I(N__13243));
    LocalMux I__1884 (
            .O(N__13243),
            .I(N__13240));
    Odrv12 I__1883 (
            .O(N__13240),
            .I(\sb_translator_1.N_1088 ));
    CEMux I__1882 (
            .O(N__13237),
            .I(N__13234));
    LocalMux I__1881 (
            .O(N__13234),
            .I(N__13231));
    Span4Mux_v I__1880 (
            .O(N__13231),
            .I(N__13228));
    Sp12to4 I__1879 (
            .O(N__13228),
            .I(N__13225));
    Odrv12 I__1878 (
            .O(N__13225),
            .I(ram_we_12));
    InMux I__1877 (
            .O(N__13222),
            .I(N__13218));
    InMux I__1876 (
            .O(N__13221),
            .I(N__13215));
    LocalMux I__1875 (
            .O(N__13218),
            .I(\spi_slave_1.mosi_data_inZ0Z_5 ));
    LocalMux I__1874 (
            .O(N__13215),
            .I(\spi_slave_1.mosi_data_inZ0Z_5 ));
    InMux I__1873 (
            .O(N__13210),
            .I(N__13206));
    InMux I__1872 (
            .O(N__13209),
            .I(N__13203));
    LocalMux I__1871 (
            .O(N__13206),
            .I(\spi_slave_1.mosi_data_inZ0Z_6 ));
    LocalMux I__1870 (
            .O(N__13203),
            .I(\spi_slave_1.mosi_data_inZ0Z_6 ));
    InMux I__1869 (
            .O(N__13198),
            .I(N__13195));
    LocalMux I__1868 (
            .O(N__13195),
            .I(N__13191));
    InMux I__1867 (
            .O(N__13194),
            .I(N__13188));
    Span4Mux_h I__1866 (
            .O(N__13191),
            .I(N__13185));
    LocalMux I__1865 (
            .O(N__13188),
            .I(\spi_slave_1.mosi_data_inZ0Z_7 ));
    Odrv4 I__1864 (
            .O(N__13185),
            .I(\spi_slave_1.mosi_data_inZ0Z_7 ));
    InMux I__1863 (
            .O(N__13180),
            .I(N__13176));
    InMux I__1862 (
            .O(N__13179),
            .I(N__13173));
    LocalMux I__1861 (
            .O(N__13176),
            .I(\spi_slave_1.mosi_data_inZ0Z_4 ));
    LocalMux I__1860 (
            .O(N__13173),
            .I(\spi_slave_1.mosi_data_inZ0Z_4 ));
    InMux I__1859 (
            .O(N__13168),
            .I(N__13164));
    InMux I__1858 (
            .O(N__13167),
            .I(N__13161));
    LocalMux I__1857 (
            .O(N__13164),
            .I(\spi_slave_1.mosi_data_inZ0Z_0 ));
    LocalMux I__1856 (
            .O(N__13161),
            .I(\spi_slave_1.mosi_data_inZ0Z_0 ));
    InMux I__1855 (
            .O(N__13156),
            .I(N__13153));
    LocalMux I__1854 (
            .O(N__13153),
            .I(N__13149));
    InMux I__1853 (
            .O(N__13152),
            .I(N__13146));
    Span4Mux_h I__1852 (
            .O(N__13149),
            .I(N__13138));
    LocalMux I__1851 (
            .O(N__13146),
            .I(N__13138));
    InMux I__1850 (
            .O(N__13145),
            .I(N__13135));
    InMux I__1849 (
            .O(N__13144),
            .I(N__13132));
    InMux I__1848 (
            .O(N__13143),
            .I(N__13129));
    Span4Mux_v I__1847 (
            .O(N__13138),
            .I(N__13120));
    LocalMux I__1846 (
            .O(N__13135),
            .I(N__13120));
    LocalMux I__1845 (
            .O(N__13132),
            .I(N__13117));
    LocalMux I__1844 (
            .O(N__13129),
            .I(N__13114));
    InMux I__1843 (
            .O(N__13128),
            .I(N__13111));
    InMux I__1842 (
            .O(N__13127),
            .I(N__13108));
    InMux I__1841 (
            .O(N__13126),
            .I(N__13104));
    InMux I__1840 (
            .O(N__13125),
            .I(N__13101));
    Span4Mux_v I__1839 (
            .O(N__13120),
            .I(N__13095));
    Span4Mux_v I__1838 (
            .O(N__13117),
            .I(N__13088));
    Span4Mux_v I__1837 (
            .O(N__13114),
            .I(N__13088));
    LocalMux I__1836 (
            .O(N__13111),
            .I(N__13088));
    LocalMux I__1835 (
            .O(N__13108),
            .I(N__13085));
    InMux I__1834 (
            .O(N__13107),
            .I(N__13082));
    LocalMux I__1833 (
            .O(N__13104),
            .I(N__13077));
    LocalMux I__1832 (
            .O(N__13101),
            .I(N__13077));
    InMux I__1831 (
            .O(N__13100),
            .I(N__13074));
    InMux I__1830 (
            .O(N__13099),
            .I(N__13071));
    InMux I__1829 (
            .O(N__13098),
            .I(N__13067));
    Span4Mux_s2_h I__1828 (
            .O(N__13095),
            .I(N__13062));
    Span4Mux_v I__1827 (
            .O(N__13088),
            .I(N__13062));
    Span4Mux_s1_v I__1826 (
            .O(N__13085),
            .I(N__13057));
    LocalMux I__1825 (
            .O(N__13082),
            .I(N__13057));
    Span4Mux_v I__1824 (
            .O(N__13077),
            .I(N__13050));
    LocalMux I__1823 (
            .O(N__13074),
            .I(N__13050));
    LocalMux I__1822 (
            .O(N__13071),
            .I(N__13050));
    InMux I__1821 (
            .O(N__13070),
            .I(N__13047));
    LocalMux I__1820 (
            .O(N__13067),
            .I(N__13044));
    Span4Mux_h I__1819 (
            .O(N__13062),
            .I(N__13035));
    Span4Mux_v I__1818 (
            .O(N__13057),
            .I(N__13035));
    Span4Mux_v I__1817 (
            .O(N__13050),
            .I(N__13035));
    LocalMux I__1816 (
            .O(N__13047),
            .I(N__13035));
    Odrv12 I__1815 (
            .O(N__13044),
            .I(ram_data_in_0));
    Odrv4 I__1814 (
            .O(N__13035),
            .I(ram_data_in_0));
    InMux I__1813 (
            .O(N__13030),
            .I(N__13025));
    InMux I__1812 (
            .O(N__13029),
            .I(N__13021));
    InMux I__1811 (
            .O(N__13028),
            .I(N__13018));
    LocalMux I__1810 (
            .O(N__13025),
            .I(N__13015));
    InMux I__1809 (
            .O(N__13024),
            .I(N__13012));
    LocalMux I__1808 (
            .O(N__13021),
            .I(N__13004));
    LocalMux I__1807 (
            .O(N__13018),
            .I(N__13001));
    Span4Mux_s1_v I__1806 (
            .O(N__13015),
            .I(N__12996));
    LocalMux I__1805 (
            .O(N__13012),
            .I(N__12996));
    InMux I__1804 (
            .O(N__13011),
            .I(N__12993));
    InMux I__1803 (
            .O(N__13010),
            .I(N__12990));
    InMux I__1802 (
            .O(N__13009),
            .I(N__12987));
    InMux I__1801 (
            .O(N__13008),
            .I(N__12983));
    InMux I__1800 (
            .O(N__13007),
            .I(N__12980));
    Span4Mux_v I__1799 (
            .O(N__13004),
            .I(N__12966));
    Span4Mux_v I__1798 (
            .O(N__13001),
            .I(N__12966));
    Span4Mux_v I__1797 (
            .O(N__12996),
            .I(N__12966));
    LocalMux I__1796 (
            .O(N__12993),
            .I(N__12966));
    LocalMux I__1795 (
            .O(N__12990),
            .I(N__12966));
    LocalMux I__1794 (
            .O(N__12987),
            .I(N__12963));
    InMux I__1793 (
            .O(N__12986),
            .I(N__12960));
    LocalMux I__1792 (
            .O(N__12983),
            .I(N__12955));
    LocalMux I__1791 (
            .O(N__12980),
            .I(N__12955));
    InMux I__1790 (
            .O(N__12979),
            .I(N__12952));
    InMux I__1789 (
            .O(N__12978),
            .I(N__12949));
    InMux I__1788 (
            .O(N__12977),
            .I(N__12945));
    Span4Mux_v I__1787 (
            .O(N__12966),
            .I(N__12942));
    Span4Mux_s1_v I__1786 (
            .O(N__12963),
            .I(N__12937));
    LocalMux I__1785 (
            .O(N__12960),
            .I(N__12937));
    Span4Mux_v I__1784 (
            .O(N__12955),
            .I(N__12930));
    LocalMux I__1783 (
            .O(N__12952),
            .I(N__12930));
    LocalMux I__1782 (
            .O(N__12949),
            .I(N__12930));
    InMux I__1781 (
            .O(N__12948),
            .I(N__12927));
    LocalMux I__1780 (
            .O(N__12945),
            .I(N__12924));
    Span4Mux_h I__1779 (
            .O(N__12942),
            .I(N__12915));
    Span4Mux_v I__1778 (
            .O(N__12937),
            .I(N__12915));
    Span4Mux_v I__1777 (
            .O(N__12930),
            .I(N__12915));
    LocalMux I__1776 (
            .O(N__12927),
            .I(N__12915));
    Odrv12 I__1775 (
            .O(N__12924),
            .I(ram_data_in_1));
    Odrv4 I__1774 (
            .O(N__12915),
            .I(ram_data_in_1));
    InMux I__1773 (
            .O(N__12910),
            .I(N__12901));
    InMux I__1772 (
            .O(N__12909),
            .I(N__12898));
    InMux I__1771 (
            .O(N__12908),
            .I(N__12891));
    InMux I__1770 (
            .O(N__12907),
            .I(N__12888));
    InMux I__1769 (
            .O(N__12906),
            .I(N__12885));
    InMux I__1768 (
            .O(N__12905),
            .I(N__12882));
    InMux I__1767 (
            .O(N__12904),
            .I(N__12879));
    LocalMux I__1766 (
            .O(N__12901),
            .I(N__12874));
    LocalMux I__1765 (
            .O(N__12898),
            .I(N__12874));
    InMux I__1764 (
            .O(N__12897),
            .I(N__12870));
    InMux I__1763 (
            .O(N__12896),
            .I(N__12867));
    InMux I__1762 (
            .O(N__12895),
            .I(N__12863));
    InMux I__1761 (
            .O(N__12894),
            .I(N__12860));
    LocalMux I__1760 (
            .O(N__12891),
            .I(N__12857));
    LocalMux I__1759 (
            .O(N__12888),
            .I(N__12851));
    LocalMux I__1758 (
            .O(N__12885),
            .I(N__12851));
    LocalMux I__1757 (
            .O(N__12882),
            .I(N__12844));
    LocalMux I__1756 (
            .O(N__12879),
            .I(N__12844));
    Span4Mux_v I__1755 (
            .O(N__12874),
            .I(N__12844));
    InMux I__1754 (
            .O(N__12873),
            .I(N__12841));
    LocalMux I__1753 (
            .O(N__12870),
            .I(N__12838));
    LocalMux I__1752 (
            .O(N__12867),
            .I(N__12835));
    InMux I__1751 (
            .O(N__12866),
            .I(N__12832));
    LocalMux I__1750 (
            .O(N__12863),
            .I(N__12829));
    LocalMux I__1749 (
            .O(N__12860),
            .I(N__12824));
    Span4Mux_h I__1748 (
            .O(N__12857),
            .I(N__12824));
    InMux I__1747 (
            .O(N__12856),
            .I(N__12821));
    Span4Mux_v I__1746 (
            .O(N__12851),
            .I(N__12816));
    Span4Mux_v I__1745 (
            .O(N__12844),
            .I(N__12816));
    LocalMux I__1744 (
            .O(N__12841),
            .I(N__12811));
    Span4Mux_s1_v I__1743 (
            .O(N__12838),
            .I(N__12811));
    Span4Mux_h I__1742 (
            .O(N__12835),
            .I(N__12808));
    LocalMux I__1741 (
            .O(N__12832),
            .I(N__12801));
    Span4Mux_h I__1740 (
            .O(N__12829),
            .I(N__12801));
    Span4Mux_v I__1739 (
            .O(N__12824),
            .I(N__12801));
    LocalMux I__1738 (
            .O(N__12821),
            .I(N__12796));
    Span4Mux_h I__1737 (
            .O(N__12816),
            .I(N__12796));
    Span4Mux_v I__1736 (
            .O(N__12811),
            .I(N__12789));
    Span4Mux_v I__1735 (
            .O(N__12808),
            .I(N__12789));
    Span4Mux_v I__1734 (
            .O(N__12801),
            .I(N__12789));
    Odrv4 I__1733 (
            .O(N__12796),
            .I(ram_data_in_2));
    Odrv4 I__1732 (
            .O(N__12789),
            .I(ram_data_in_2));
    InMux I__1731 (
            .O(N__12784),
            .I(N__12780));
    InMux I__1730 (
            .O(N__12783),
            .I(N__12772));
    LocalMux I__1729 (
            .O(N__12780),
            .I(N__12768));
    InMux I__1728 (
            .O(N__12779),
            .I(N__12765));
    InMux I__1727 (
            .O(N__12778),
            .I(N__12762));
    InMux I__1726 (
            .O(N__12777),
            .I(N__12758));
    InMux I__1725 (
            .O(N__12776),
            .I(N__12754));
    InMux I__1724 (
            .O(N__12775),
            .I(N__12748));
    LocalMux I__1723 (
            .O(N__12772),
            .I(N__12745));
    InMux I__1722 (
            .O(N__12771),
            .I(N__12742));
    Span4Mux_h I__1721 (
            .O(N__12768),
            .I(N__12737));
    LocalMux I__1720 (
            .O(N__12765),
            .I(N__12737));
    LocalMux I__1719 (
            .O(N__12762),
            .I(N__12734));
    InMux I__1718 (
            .O(N__12761),
            .I(N__12731));
    LocalMux I__1717 (
            .O(N__12758),
            .I(N__12728));
    InMux I__1716 (
            .O(N__12757),
            .I(N__12725));
    LocalMux I__1715 (
            .O(N__12754),
            .I(N__12722));
    InMux I__1714 (
            .O(N__12753),
            .I(N__12719));
    InMux I__1713 (
            .O(N__12752),
            .I(N__12716));
    InMux I__1712 (
            .O(N__12751),
            .I(N__12713));
    LocalMux I__1711 (
            .O(N__12748),
            .I(N__12710));
    Span4Mux_s1_v I__1710 (
            .O(N__12745),
            .I(N__12705));
    LocalMux I__1709 (
            .O(N__12742),
            .I(N__12705));
    Span4Mux_v I__1708 (
            .O(N__12737),
            .I(N__12698));
    Span4Mux_h I__1707 (
            .O(N__12734),
            .I(N__12698));
    LocalMux I__1706 (
            .O(N__12731),
            .I(N__12698));
    Span4Mux_s1_v I__1705 (
            .O(N__12728),
            .I(N__12693));
    LocalMux I__1704 (
            .O(N__12725),
            .I(N__12693));
    Sp12to4 I__1703 (
            .O(N__12722),
            .I(N__12683));
    LocalMux I__1702 (
            .O(N__12719),
            .I(N__12683));
    LocalMux I__1701 (
            .O(N__12716),
            .I(N__12683));
    LocalMux I__1700 (
            .O(N__12713),
            .I(N__12683));
    Span4Mux_h I__1699 (
            .O(N__12710),
            .I(N__12676));
    Span4Mux_v I__1698 (
            .O(N__12705),
            .I(N__12676));
    Span4Mux_v I__1697 (
            .O(N__12698),
            .I(N__12676));
    Span4Mux_v I__1696 (
            .O(N__12693),
            .I(N__12673));
    InMux I__1695 (
            .O(N__12692),
            .I(N__12670));
    Span12Mux_s8_v I__1694 (
            .O(N__12683),
            .I(N__12665));
    Sp12to4 I__1693 (
            .O(N__12676),
            .I(N__12665));
    Span4Mux_h I__1692 (
            .O(N__12673),
            .I(N__12660));
    LocalMux I__1691 (
            .O(N__12670),
            .I(N__12660));
    Odrv12 I__1690 (
            .O(N__12665),
            .I(ram_data_in_3));
    Odrv4 I__1689 (
            .O(N__12660),
            .I(ram_data_in_3));
    InMux I__1688 (
            .O(N__12655),
            .I(N__12647));
    InMux I__1687 (
            .O(N__12654),
            .I(N__12644));
    InMux I__1686 (
            .O(N__12653),
            .I(N__12637));
    InMux I__1685 (
            .O(N__12652),
            .I(N__12632));
    InMux I__1684 (
            .O(N__12651),
            .I(N__12627));
    InMux I__1683 (
            .O(N__12650),
            .I(N__12624));
    LocalMux I__1682 (
            .O(N__12647),
            .I(N__12619));
    LocalMux I__1681 (
            .O(N__12644),
            .I(N__12619));
    InMux I__1680 (
            .O(N__12643),
            .I(N__12616));
    InMux I__1679 (
            .O(N__12642),
            .I(N__12613));
    InMux I__1678 (
            .O(N__12641),
            .I(N__12610));
    InMux I__1677 (
            .O(N__12640),
            .I(N__12607));
    LocalMux I__1676 (
            .O(N__12637),
            .I(N__12604));
    InMux I__1675 (
            .O(N__12636),
            .I(N__12601));
    InMux I__1674 (
            .O(N__12635),
            .I(N__12598));
    LocalMux I__1673 (
            .O(N__12632),
            .I(N__12595));
    InMux I__1672 (
            .O(N__12631),
            .I(N__12592));
    InMux I__1671 (
            .O(N__12630),
            .I(N__12589));
    LocalMux I__1670 (
            .O(N__12627),
            .I(N__12584));
    LocalMux I__1669 (
            .O(N__12624),
            .I(N__12584));
    Span4Mux_s3_v I__1668 (
            .O(N__12619),
            .I(N__12577));
    LocalMux I__1667 (
            .O(N__12616),
            .I(N__12577));
    LocalMux I__1666 (
            .O(N__12613),
            .I(N__12577));
    LocalMux I__1665 (
            .O(N__12610),
            .I(N__12574));
    LocalMux I__1664 (
            .O(N__12607),
            .I(N__12569));
    Span4Mux_s2_v I__1663 (
            .O(N__12604),
            .I(N__12569));
    LocalMux I__1662 (
            .O(N__12601),
            .I(N__12566));
    LocalMux I__1661 (
            .O(N__12598),
            .I(N__12561));
    Span4Mux_s1_v I__1660 (
            .O(N__12595),
            .I(N__12561));
    LocalMux I__1659 (
            .O(N__12592),
            .I(N__12554));
    LocalMux I__1658 (
            .O(N__12589),
            .I(N__12554));
    Span4Mux_v I__1657 (
            .O(N__12584),
            .I(N__12554));
    Span4Mux_v I__1656 (
            .O(N__12577),
            .I(N__12547));
    Span4Mux_v I__1655 (
            .O(N__12574),
            .I(N__12547));
    Span4Mux_v I__1654 (
            .O(N__12569),
            .I(N__12547));
    Span4Mux_v I__1653 (
            .O(N__12566),
            .I(N__12540));
    Span4Mux_v I__1652 (
            .O(N__12561),
            .I(N__12540));
    Span4Mux_v I__1651 (
            .O(N__12554),
            .I(N__12540));
    Span4Mux_h I__1650 (
            .O(N__12547),
            .I(N__12537));
    Odrv4 I__1649 (
            .O(N__12540),
            .I(ram_data_in_4));
    Odrv4 I__1648 (
            .O(N__12537),
            .I(ram_data_in_4));
    InMux I__1647 (
            .O(N__12532),
            .I(N__12526));
    InMux I__1646 (
            .O(N__12531),
            .I(N__12526));
    LocalMux I__1645 (
            .O(N__12526),
            .I(N__12523));
    Span4Mux_h I__1644 (
            .O(N__12523),
            .I(N__12520));
    Odrv4 I__1643 (
            .O(N__12520),
            .I(mosi_data_out_8));
    InMux I__1642 (
            .O(N__12517),
            .I(N__12514));
    LocalMux I__1641 (
            .O(N__12514),
            .I(N__12509));
    InMux I__1640 (
            .O(N__12513),
            .I(N__12505));
    InMux I__1639 (
            .O(N__12512),
            .I(N__12502));
    Span4Mux_v I__1638 (
            .O(N__12509),
            .I(N__12499));
    InMux I__1637 (
            .O(N__12508),
            .I(N__12496));
    LocalMux I__1636 (
            .O(N__12505),
            .I(N__12493));
    LocalMux I__1635 (
            .O(N__12502),
            .I(\sb_translator_1.cntZ0Z_0 ));
    Odrv4 I__1634 (
            .O(N__12499),
            .I(\sb_translator_1.cntZ0Z_0 ));
    LocalMux I__1633 (
            .O(N__12496),
            .I(\sb_translator_1.cntZ0Z_0 ));
    Odrv4 I__1632 (
            .O(N__12493),
            .I(\sb_translator_1.cntZ0Z_0 ));
    InMux I__1631 (
            .O(N__12484),
            .I(N__12478));
    InMux I__1630 (
            .O(N__12483),
            .I(N__12478));
    LocalMux I__1629 (
            .O(N__12478),
            .I(N__12475));
    Odrv4 I__1628 (
            .O(N__12475),
            .I(mosi_data_out_9));
    InMux I__1627 (
            .O(N__12472),
            .I(N__12468));
    InMux I__1626 (
            .O(N__12471),
            .I(N__12465));
    LocalMux I__1625 (
            .O(N__12468),
            .I(N__12462));
    LocalMux I__1624 (
            .O(N__12465),
            .I(N__12458));
    Span4Mux_h I__1623 (
            .O(N__12462),
            .I(N__12455));
    InMux I__1622 (
            .O(N__12461),
            .I(N__12452));
    Span4Mux_s2_h I__1621 (
            .O(N__12458),
            .I(N__12449));
    Odrv4 I__1620 (
            .O(N__12455),
            .I(\sb_translator_1.cntZ0Z_1 ));
    LocalMux I__1619 (
            .O(N__12452),
            .I(\sb_translator_1.cntZ0Z_1 ));
    Odrv4 I__1618 (
            .O(N__12449),
            .I(\sb_translator_1.cntZ0Z_1 ));
    InMux I__1617 (
            .O(N__12442),
            .I(N__12439));
    LocalMux I__1616 (
            .O(N__12439),
            .I(N__12435));
    InMux I__1615 (
            .O(N__12438),
            .I(N__12431));
    Span4Mux_v I__1614 (
            .O(N__12435),
            .I(N__12428));
    InMux I__1613 (
            .O(N__12434),
            .I(N__12425));
    LocalMux I__1612 (
            .O(N__12431),
            .I(N__12422));
    Odrv4 I__1611 (
            .O(N__12428),
            .I(\sb_translator_1.cntZ0Z_2 ));
    LocalMux I__1610 (
            .O(N__12425),
            .I(\sb_translator_1.cntZ0Z_2 ));
    Odrv4 I__1609 (
            .O(N__12422),
            .I(\sb_translator_1.cntZ0Z_2 ));
    InMux I__1608 (
            .O(N__12415),
            .I(N__12409));
    InMux I__1607 (
            .O(N__12414),
            .I(N__12409));
    LocalMux I__1606 (
            .O(N__12409),
            .I(N__12406));
    Odrv12 I__1605 (
            .O(N__12406),
            .I(mosi_data_out_10));
    InMux I__1604 (
            .O(N__12403),
            .I(N__12400));
    LocalMux I__1603 (
            .O(N__12400),
            .I(N__12396));
    InMux I__1602 (
            .O(N__12399),
            .I(N__12393));
    Odrv12 I__1601 (
            .O(N__12396),
            .I(\spi_slave_1.mosi_data_inZ0Z_16 ));
    LocalMux I__1600 (
            .O(N__12393),
            .I(\spi_slave_1.mosi_data_inZ0Z_16 ));
    InMux I__1599 (
            .O(N__12388),
            .I(N__12384));
    InMux I__1598 (
            .O(N__12387),
            .I(N__12381));
    LocalMux I__1597 (
            .O(N__12384),
            .I(\spi_slave_1.mosi_data_inZ0Z_3 ));
    LocalMux I__1596 (
            .O(N__12381),
            .I(\spi_slave_1.mosi_data_inZ0Z_3 ));
    InMux I__1595 (
            .O(N__12376),
            .I(N__12372));
    InMux I__1594 (
            .O(N__12375),
            .I(N__12369));
    LocalMux I__1593 (
            .O(N__12372),
            .I(\spi_slave_1.mosi_data_inZ0Z_2 ));
    LocalMux I__1592 (
            .O(N__12369),
            .I(\spi_slave_1.mosi_data_inZ0Z_2 ));
    InMux I__1591 (
            .O(N__12364),
            .I(N__12331));
    InMux I__1590 (
            .O(N__12363),
            .I(N__12331));
    InMux I__1589 (
            .O(N__12362),
            .I(N__12331));
    InMux I__1588 (
            .O(N__12361),
            .I(N__12331));
    InMux I__1587 (
            .O(N__12360),
            .I(N__12331));
    InMux I__1586 (
            .O(N__12359),
            .I(N__12331));
    InMux I__1585 (
            .O(N__12358),
            .I(N__12331));
    InMux I__1584 (
            .O(N__12357),
            .I(N__12331));
    InMux I__1583 (
            .O(N__12356),
            .I(N__12306));
    InMux I__1582 (
            .O(N__12355),
            .I(N__12306));
    InMux I__1581 (
            .O(N__12354),
            .I(N__12306));
    InMux I__1580 (
            .O(N__12353),
            .I(N__12306));
    InMux I__1579 (
            .O(N__12352),
            .I(N__12306));
    InMux I__1578 (
            .O(N__12351),
            .I(N__12306));
    InMux I__1577 (
            .O(N__12350),
            .I(N__12306));
    InMux I__1576 (
            .O(N__12349),
            .I(N__12306));
    InMux I__1575 (
            .O(N__12348),
            .I(N__12303));
    LocalMux I__1574 (
            .O(N__12331),
            .I(N__12300));
    InMux I__1573 (
            .O(N__12330),
            .I(N__12283));
    InMux I__1572 (
            .O(N__12329),
            .I(N__12283));
    InMux I__1571 (
            .O(N__12328),
            .I(N__12283));
    InMux I__1570 (
            .O(N__12327),
            .I(N__12283));
    InMux I__1569 (
            .O(N__12326),
            .I(N__12283));
    InMux I__1568 (
            .O(N__12325),
            .I(N__12283));
    InMux I__1567 (
            .O(N__12324),
            .I(N__12283));
    InMux I__1566 (
            .O(N__12323),
            .I(N__12283));
    LocalMux I__1565 (
            .O(N__12306),
            .I(N__12278));
    LocalMux I__1564 (
            .O(N__12303),
            .I(N__12278));
    Span4Mux_h I__1563 (
            .O(N__12300),
            .I(N__12270));
    LocalMux I__1562 (
            .O(N__12283),
            .I(N__12270));
    Span4Mux_h I__1561 (
            .O(N__12278),
            .I(N__12270));
    InMux I__1560 (
            .O(N__12277),
            .I(N__12264));
    Sp12to4 I__1559 (
            .O(N__12270),
            .I(N__12261));
    InMux I__1558 (
            .O(N__12269),
            .I(N__12254));
    InMux I__1557 (
            .O(N__12268),
            .I(N__12254));
    InMux I__1556 (
            .O(N__12267),
            .I(N__12254));
    LocalMux I__1555 (
            .O(N__12264),
            .I(\spi_slave_1.clkZ0Z_0 ));
    Odrv12 I__1554 (
            .O(N__12261),
            .I(\spi_slave_1.clkZ0Z_0 ));
    LocalMux I__1553 (
            .O(N__12254),
            .I(\spi_slave_1.clkZ0Z_0 ));
    CascadeMux I__1552 (
            .O(N__12247),
            .I(N__12241));
    CascadeMux I__1551 (
            .O(N__12246),
            .I(N__12237));
    CascadeMux I__1550 (
            .O(N__12245),
            .I(N__12233));
    CascadeMux I__1549 (
            .O(N__12244),
            .I(N__12229));
    InMux I__1548 (
            .O(N__12241),
            .I(N__12203));
    InMux I__1547 (
            .O(N__12240),
            .I(N__12203));
    InMux I__1546 (
            .O(N__12237),
            .I(N__12203));
    InMux I__1545 (
            .O(N__12236),
            .I(N__12203));
    InMux I__1544 (
            .O(N__12233),
            .I(N__12203));
    InMux I__1543 (
            .O(N__12232),
            .I(N__12203));
    InMux I__1542 (
            .O(N__12229),
            .I(N__12203));
    InMux I__1541 (
            .O(N__12228),
            .I(N__12203));
    CascadeMux I__1540 (
            .O(N__12227),
            .I(N__12199));
    CascadeMux I__1539 (
            .O(N__12226),
            .I(N__12195));
    CascadeMux I__1538 (
            .O(N__12225),
            .I(N__12191));
    CascadeMux I__1537 (
            .O(N__12224),
            .I(N__12187));
    CascadeMux I__1536 (
            .O(N__12223),
            .I(N__12183));
    CascadeMux I__1535 (
            .O(N__12222),
            .I(N__12179));
    CascadeMux I__1534 (
            .O(N__12221),
            .I(N__12175));
    CascadeMux I__1533 (
            .O(N__12220),
            .I(N__12171));
    LocalMux I__1532 (
            .O(N__12203),
            .I(N__12167));
    InMux I__1531 (
            .O(N__12202),
            .I(N__12164));
    InMux I__1530 (
            .O(N__12199),
            .I(N__12147));
    InMux I__1529 (
            .O(N__12198),
            .I(N__12147));
    InMux I__1528 (
            .O(N__12195),
            .I(N__12147));
    InMux I__1527 (
            .O(N__12194),
            .I(N__12147));
    InMux I__1526 (
            .O(N__12191),
            .I(N__12147));
    InMux I__1525 (
            .O(N__12190),
            .I(N__12147));
    InMux I__1524 (
            .O(N__12187),
            .I(N__12147));
    InMux I__1523 (
            .O(N__12186),
            .I(N__12147));
    InMux I__1522 (
            .O(N__12183),
            .I(N__12129));
    InMux I__1521 (
            .O(N__12182),
            .I(N__12129));
    InMux I__1520 (
            .O(N__12179),
            .I(N__12129));
    InMux I__1519 (
            .O(N__12178),
            .I(N__12129));
    InMux I__1518 (
            .O(N__12175),
            .I(N__12129));
    InMux I__1517 (
            .O(N__12174),
            .I(N__12129));
    InMux I__1516 (
            .O(N__12171),
            .I(N__12129));
    InMux I__1515 (
            .O(N__12170),
            .I(N__12129));
    Span4Mux_v I__1514 (
            .O(N__12167),
            .I(N__12124));
    LocalMux I__1513 (
            .O(N__12164),
            .I(N__12124));
    LocalMux I__1512 (
            .O(N__12147),
            .I(N__12121));
    InMux I__1511 (
            .O(N__12146),
            .I(N__12118));
    LocalMux I__1510 (
            .O(N__12129),
            .I(N__12113));
    Sp12to4 I__1509 (
            .O(N__12124),
            .I(N__12113));
    Span12Mux_s3_v I__1508 (
            .O(N__12121),
            .I(N__12108));
    LocalMux I__1507 (
            .O(N__12118),
            .I(N__12105));
    Span12Mux_s10_v I__1506 (
            .O(N__12113),
            .I(N__12102));
    InMux I__1505 (
            .O(N__12112),
            .I(N__12097));
    InMux I__1504 (
            .O(N__12111),
            .I(N__12097));
    Odrv12 I__1503 (
            .O(N__12108),
            .I(\spi_slave_1.clkZ0Z_1 ));
    Odrv4 I__1502 (
            .O(N__12105),
            .I(\spi_slave_1.clkZ0Z_1 ));
    Odrv12 I__1501 (
            .O(N__12102),
            .I(\spi_slave_1.clkZ0Z_1 ));
    LocalMux I__1500 (
            .O(N__12097),
            .I(\spi_slave_1.clkZ0Z_1 ));
    InMux I__1499 (
            .O(N__12088),
            .I(N__12084));
    InMux I__1498 (
            .O(N__12087),
            .I(N__12081));
    LocalMux I__1497 (
            .O(N__12084),
            .I(N__12078));
    LocalMux I__1496 (
            .O(N__12081),
            .I(N__12075));
    Span4Mux_h I__1495 (
            .O(N__12078),
            .I(N__12072));
    Span4Mux_h I__1494 (
            .O(N__12075),
            .I(N__12069));
    Odrv4 I__1493 (
            .O(N__12072),
            .I(\spi_slave_1.mosi_data_inZ0Z_17 ));
    Odrv4 I__1492 (
            .O(N__12069),
            .I(\spi_slave_1.mosi_data_inZ0Z_17 ));
    CEMux I__1491 (
            .O(N__12064),
            .I(N__12052));
    CEMux I__1490 (
            .O(N__12063),
            .I(N__12052));
    CEMux I__1489 (
            .O(N__12062),
            .I(N__12052));
    CEMux I__1488 (
            .O(N__12061),
            .I(N__12052));
    GlobalMux I__1487 (
            .O(N__12052),
            .I(N__12049));
    gio2CtrlBuf I__1486 (
            .O(N__12049),
            .I(\spi_slave_1.bitcnt_rxe_0_i_g ));
    InMux I__1485 (
            .O(N__12046),
            .I(N__12042));
    InMux I__1484 (
            .O(N__12045),
            .I(N__12039));
    LocalMux I__1483 (
            .O(N__12042),
            .I(N__12036));
    LocalMux I__1482 (
            .O(N__12039),
            .I(N__12033));
    Span4Mux_h I__1481 (
            .O(N__12036),
            .I(N__12030));
    Span4Mux_h I__1480 (
            .O(N__12033),
            .I(N__12027));
    Odrv4 I__1479 (
            .O(N__12030),
            .I(\spi_slave_1.mosi_data_inZ0Z_9 ));
    Odrv4 I__1478 (
            .O(N__12027),
            .I(\spi_slave_1.mosi_data_inZ0Z_9 ));
    InMux I__1477 (
            .O(N__12022),
            .I(N__12019));
    LocalMux I__1476 (
            .O(N__12019),
            .I(N__12016));
    Span4Mux_h I__1475 (
            .O(N__12016),
            .I(N__12012));
    InMux I__1474 (
            .O(N__12015),
            .I(N__12009));
    Odrv4 I__1473 (
            .O(N__12012),
            .I(\spi_slave_1.mosi_data_inZ0Z_8 ));
    LocalMux I__1472 (
            .O(N__12009),
            .I(\spi_slave_1.mosi_data_inZ0Z_8 ));
    InMux I__1471 (
            .O(N__12004),
            .I(N__12000));
    InMux I__1470 (
            .O(N__12003),
            .I(N__11997));
    LocalMux I__1469 (
            .O(N__12000),
            .I(\spi_slave_1.mosi_data_inZ0Z_10 ));
    LocalMux I__1468 (
            .O(N__11997),
            .I(\spi_slave_1.mosi_data_inZ0Z_10 ));
    InMux I__1467 (
            .O(N__11992),
            .I(N__11988));
    InMux I__1466 (
            .O(N__11991),
            .I(N__11985));
    LocalMux I__1465 (
            .O(N__11988),
            .I(\spi_slave_1.mosi_data_inZ0Z_11 ));
    LocalMux I__1464 (
            .O(N__11985),
            .I(\spi_slave_1.mosi_data_inZ0Z_11 ));
    InMux I__1463 (
            .O(N__11980),
            .I(N__11976));
    InMux I__1462 (
            .O(N__11979),
            .I(N__11973));
    LocalMux I__1461 (
            .O(N__11976),
            .I(\spi_slave_1.mosi_data_inZ0Z_12 ));
    LocalMux I__1460 (
            .O(N__11973),
            .I(\spi_slave_1.mosi_data_inZ0Z_12 ));
    InMux I__1459 (
            .O(N__11968),
            .I(N__11964));
    InMux I__1458 (
            .O(N__11967),
            .I(N__11961));
    LocalMux I__1457 (
            .O(N__11964),
            .I(\spi_slave_1.mosi_data_inZ0Z_13 ));
    LocalMux I__1456 (
            .O(N__11961),
            .I(\spi_slave_1.mosi_data_inZ0Z_13 ));
    InMux I__1455 (
            .O(N__11956),
            .I(N__11952));
    InMux I__1454 (
            .O(N__11955),
            .I(N__11949));
    LocalMux I__1453 (
            .O(N__11952),
            .I(\spi_slave_1.mosi_data_inZ0Z_14 ));
    LocalMux I__1452 (
            .O(N__11949),
            .I(\spi_slave_1.mosi_data_inZ0Z_14 ));
    InMux I__1451 (
            .O(N__11944),
            .I(N__11936));
    InMux I__1450 (
            .O(N__11943),
            .I(N__11936));
    InMux I__1449 (
            .O(N__11942),
            .I(N__11928));
    InMux I__1448 (
            .O(N__11941),
            .I(N__11928));
    LocalMux I__1447 (
            .O(N__11936),
            .I(N__11925));
    InMux I__1446 (
            .O(N__11935),
            .I(N__11918));
    InMux I__1445 (
            .O(N__11934),
            .I(N__11918));
    InMux I__1444 (
            .O(N__11933),
            .I(N__11918));
    LocalMux I__1443 (
            .O(N__11928),
            .I(\spi_slave_1.bitcnt_txZ0Z_1 ));
    Odrv12 I__1442 (
            .O(N__11925),
            .I(\spi_slave_1.bitcnt_txZ0Z_1 ));
    LocalMux I__1441 (
            .O(N__11918),
            .I(\spi_slave_1.bitcnt_txZ0Z_1 ));
    CascadeMux I__1440 (
            .O(N__11911),
            .I(\spi_slave_1.m27_ns_1_cascade_ ));
    InMux I__1439 (
            .O(N__11908),
            .I(N__11905));
    LocalMux I__1438 (
            .O(N__11905),
            .I(N__11902));
    Span4Mux_s3_v I__1437 (
            .O(N__11902),
            .I(N__11899));
    Odrv4 I__1436 (
            .O(N__11899),
            .I(\spi_slave_1.miso_RNOZ0Z_7 ));
    InMux I__1435 (
            .O(N__11896),
            .I(N__11893));
    LocalMux I__1434 (
            .O(N__11893),
            .I(N__11890));
    Odrv4 I__1433 (
            .O(N__11890),
            .I(\spi_slave_1.N_28_0 ));
    InMux I__1432 (
            .O(N__11887),
            .I(N__11884));
    LocalMux I__1431 (
            .O(N__11884),
            .I(N__11881));
    Odrv12 I__1430 (
            .O(N__11881),
            .I(\spi_slave_1.mosi_bufferZ0Z_1 ));
    InMux I__1429 (
            .O(N__11878),
            .I(N__11873));
    CascadeMux I__1428 (
            .O(N__11877),
            .I(N__11870));
    CascadeMux I__1427 (
            .O(N__11876),
            .I(N__11865));
    LocalMux I__1426 (
            .O(N__11873),
            .I(N__11859));
    InMux I__1425 (
            .O(N__11870),
            .I(N__11856));
    InMux I__1424 (
            .O(N__11869),
            .I(N__11851));
    InMux I__1423 (
            .O(N__11868),
            .I(N__11851));
    InMux I__1422 (
            .O(N__11865),
            .I(N__11848));
    CascadeMux I__1421 (
            .O(N__11864),
            .I(N__11845));
    CascadeMux I__1420 (
            .O(N__11863),
            .I(N__11842));
    CascadeMux I__1419 (
            .O(N__11862),
            .I(N__11838));
    Span12Mux_s11_h I__1418 (
            .O(N__11859),
            .I(N__11835));
    LocalMux I__1417 (
            .O(N__11856),
            .I(N__11832));
    LocalMux I__1416 (
            .O(N__11851),
            .I(N__11829));
    LocalMux I__1415 (
            .O(N__11848),
            .I(N__11826));
    InMux I__1414 (
            .O(N__11845),
            .I(N__11823));
    InMux I__1413 (
            .O(N__11842),
            .I(N__11820));
    InMux I__1412 (
            .O(N__11841),
            .I(N__11815));
    InMux I__1411 (
            .O(N__11838),
            .I(N__11815));
    Span12Mux_v I__1410 (
            .O(N__11835),
            .I(N__11812));
    Span4Mux_v I__1409 (
            .O(N__11832),
            .I(N__11807));
    Span4Mux_h I__1408 (
            .O(N__11829),
            .I(N__11807));
    Span12Mux_s2_h I__1407 (
            .O(N__11826),
            .I(N__11798));
    LocalMux I__1406 (
            .O(N__11823),
            .I(N__11798));
    LocalMux I__1405 (
            .O(N__11820),
            .I(N__11798));
    LocalMux I__1404 (
            .O(N__11815),
            .I(N__11798));
    Odrv12 I__1403 (
            .O(N__11812),
            .I(cs_n));
    Odrv4 I__1402 (
            .O(N__11807),
            .I(cs_n));
    Odrv12 I__1401 (
            .O(N__11798),
            .I(cs_n));
    InMux I__1400 (
            .O(N__11791),
            .I(N__11788));
    LocalMux I__1399 (
            .O(N__11788),
            .I(N__11785));
    IoSpan4Mux I__1398 (
            .O(N__11785),
            .I(N__11782));
    IoSpan4Mux I__1397 (
            .O(N__11782),
            .I(N__11779));
    Odrv4 I__1396 (
            .O(N__11779),
            .I(mosi));
    InMux I__1395 (
            .O(N__11776),
            .I(N__11773));
    LocalMux I__1394 (
            .O(N__11773),
            .I(\spi_slave_1.mosi_bufferZ0Z_0 ));
    InMux I__1393 (
            .O(N__11770),
            .I(N__11767));
    LocalMux I__1392 (
            .O(N__11767),
            .I(N__11764));
    Span4Mux_h I__1391 (
            .O(N__11764),
            .I(N__11761));
    Odrv4 I__1390 (
            .O(N__11761),
            .I(\spi_slave_1.miso_data_outZ0Z_3 ));
    InMux I__1389 (
            .O(N__11758),
            .I(N__11755));
    LocalMux I__1388 (
            .O(N__11755),
            .I(N__11752));
    Odrv4 I__1387 (
            .O(N__11752),
            .I(\spi_slave_1.miso_data_outZ0Z_7 ));
    InMux I__1386 (
            .O(N__11749),
            .I(N__11746));
    LocalMux I__1385 (
            .O(N__11746),
            .I(N__11743));
    Span4Mux_v I__1384 (
            .O(N__11743),
            .I(N__11740));
    Odrv4 I__1383 (
            .O(N__11740),
            .I(miso_data_in_18));
    InMux I__1382 (
            .O(N__11737),
            .I(N__11734));
    LocalMux I__1381 (
            .O(N__11734),
            .I(\spi_slave_1.miso_data_outZ0Z_2 ));
    CascadeMux I__1380 (
            .O(N__11731),
            .I(N__11728));
    InMux I__1379 (
            .O(N__11728),
            .I(N__11725));
    LocalMux I__1378 (
            .O(N__11725),
            .I(\spi_slave_1.miso_data_outZ0Z_18 ));
    InMux I__1377 (
            .O(N__11722),
            .I(N__11719));
    LocalMux I__1376 (
            .O(N__11719),
            .I(N__11716));
    Span4Mux_v I__1375 (
            .O(N__11716),
            .I(N__11713));
    Odrv4 I__1374 (
            .O(N__11713),
            .I(\spi_slave_1.m72_ns_1 ));
    InMux I__1373 (
            .O(N__11710),
            .I(N__11707));
    LocalMux I__1372 (
            .O(N__11707),
            .I(\spi_slave_1.miso_data_outZ0Z_14 ));
    InMux I__1371 (
            .O(N__11704),
            .I(N__11701));
    LocalMux I__1370 (
            .O(N__11701),
            .I(\spi_slave_1.miso_data_outZ0Z_13 ));
    InMux I__1369 (
            .O(N__11698),
            .I(N__11691));
    CascadeMux I__1368 (
            .O(N__11697),
            .I(N__11688));
    CascadeMux I__1367 (
            .O(N__11696),
            .I(N__11685));
    InMux I__1366 (
            .O(N__11695),
            .I(N__11680));
    InMux I__1365 (
            .O(N__11694),
            .I(N__11680));
    LocalMux I__1364 (
            .O(N__11691),
            .I(N__11677));
    InMux I__1363 (
            .O(N__11688),
            .I(N__11672));
    InMux I__1362 (
            .O(N__11685),
            .I(N__11672));
    LocalMux I__1361 (
            .O(N__11680),
            .I(\spi_slave_1.bitcnt_txZ0Z_2 ));
    Odrv4 I__1360 (
            .O(N__11677),
            .I(\spi_slave_1.bitcnt_txZ0Z_2 ));
    LocalMux I__1359 (
            .O(N__11672),
            .I(\spi_slave_1.bitcnt_txZ0Z_2 ));
    CascadeMux I__1358 (
            .O(N__11665),
            .I(\spi_slave_1.miso_RNOZ0Z_12_cascade_ ));
    InMux I__1357 (
            .O(N__11662),
            .I(N__11659));
    LocalMux I__1356 (
            .O(N__11659),
            .I(N__11656));
    Span4Mux_v I__1355 (
            .O(N__11656),
            .I(N__11653));
    Odrv4 I__1354 (
            .O(N__11653),
            .I(demux_data_in_55));
    CascadeMux I__1353 (
            .O(N__11650),
            .I(\demux.N_417_i_0_o2Z0Z_6_cascade_ ));
    InMux I__1352 (
            .O(N__11647),
            .I(N__11644));
    LocalMux I__1351 (
            .O(N__11644),
            .I(\demux.N_890 ));
    InMux I__1350 (
            .O(N__11641),
            .I(N__11638));
    LocalMux I__1349 (
            .O(N__11638),
            .I(demux_data_in_61));
    InMux I__1348 (
            .O(N__11635),
            .I(N__11632));
    LocalMux I__1347 (
            .O(N__11632),
            .I(N__11629));
    Span4Mux_v I__1346 (
            .O(N__11629),
            .I(N__11626));
    Odrv4 I__1345 (
            .O(N__11626),
            .I(demux_data_in_77));
    CascadeMux I__1344 (
            .O(N__11623),
            .I(N__11620));
    InMux I__1343 (
            .O(N__11620),
            .I(N__11617));
    LocalMux I__1342 (
            .O(N__11617),
            .I(N__11614));
    Span4Mux_h I__1341 (
            .O(N__11614),
            .I(N__11611));
    Span4Mux_h I__1340 (
            .O(N__11611),
            .I(N__11608));
    Span4Mux_v I__1339 (
            .O(N__11608),
            .I(N__11605));
    Odrv4 I__1338 (
            .O(N__11605),
            .I(demux_data_in_85));
    InMux I__1337 (
            .O(N__11602),
            .I(N__11599));
    LocalMux I__1336 (
            .O(N__11599),
            .I(N__11596));
    Span4Mux_h I__1335 (
            .O(N__11596),
            .I(N__11593));
    Span4Mux_s3_h I__1334 (
            .O(N__11593),
            .I(N__11590));
    Odrv4 I__1333 (
            .O(N__11590),
            .I(demux_data_in_53));
    CascadeMux I__1332 (
            .O(N__11587),
            .I(\demux.N_419_i_0_o2Z0Z_6_cascade_ ));
    InMux I__1331 (
            .O(N__11584),
            .I(N__11581));
    LocalMux I__1330 (
            .O(N__11581),
            .I(\demux.N_419_i_0_a3Z0Z_1 ));
    InMux I__1329 (
            .O(N__11578),
            .I(N__11575));
    LocalMux I__1328 (
            .O(N__11575),
            .I(demux_data_in_60));
    InMux I__1327 (
            .O(N__11572),
            .I(N__11569));
    LocalMux I__1326 (
            .O(N__11569),
            .I(N__11566));
    Span4Mux_h I__1325 (
            .O(N__11566),
            .I(N__11563));
    Span4Mux_h I__1324 (
            .O(N__11563),
            .I(N__11560));
    Span4Mux_v I__1323 (
            .O(N__11560),
            .I(N__11557));
    Odrv4 I__1322 (
            .O(N__11557),
            .I(demux_data_in_84));
    InMux I__1321 (
            .O(N__11554),
            .I(N__11551));
    LocalMux I__1320 (
            .O(N__11551),
            .I(N__11548));
    Span4Mux_h I__1319 (
            .O(N__11548),
            .I(N__11545));
    Odrv4 I__1318 (
            .O(N__11545),
            .I(demux_data_in_76));
    InMux I__1317 (
            .O(N__11542),
            .I(N__11539));
    LocalMux I__1316 (
            .O(N__11539),
            .I(N__11536));
    Odrv4 I__1315 (
            .O(N__11536),
            .I(demux_data_in_52));
    CascadeMux I__1314 (
            .O(N__11533),
            .I(\demux.N_420_i_0_o2Z0Z_6_cascade_ ));
    InMux I__1313 (
            .O(N__11530),
            .I(N__11527));
    LocalMux I__1312 (
            .O(N__11527),
            .I(\demux.N_420_i_0_a3Z0Z_1 ));
    InMux I__1311 (
            .O(N__11524),
            .I(N__11521));
    LocalMux I__1310 (
            .O(N__11521),
            .I(N__11518));
    Span4Mux_v I__1309 (
            .O(N__11518),
            .I(N__11515));
    Odrv4 I__1308 (
            .O(N__11515),
            .I(\spi_slave_1.miso_data_outZ0Z_6 ));
    InMux I__1307 (
            .O(N__11512),
            .I(N__11509));
    LocalMux I__1306 (
            .O(N__11509),
            .I(N__11506));
    Odrv4 I__1305 (
            .O(N__11506),
            .I(\spi_slave_1.miso_data_outZ0Z_1 ));
    InMux I__1304 (
            .O(N__11503),
            .I(N__11500));
    LocalMux I__1303 (
            .O(N__11500),
            .I(N__11497));
    Odrv4 I__1302 (
            .O(N__11497),
            .I(demux_data_in_54));
    CascadeMux I__1301 (
            .O(N__11494),
            .I(\demux.N_877_cascade_ ));
    InMux I__1300 (
            .O(N__11491),
            .I(N__11488));
    LocalMux I__1299 (
            .O(N__11488),
            .I(N__11485));
    Odrv4 I__1298 (
            .O(N__11485),
            .I(demux_data_in_70));
    InMux I__1297 (
            .O(N__11482),
            .I(N__11479));
    LocalMux I__1296 (
            .O(N__11479),
            .I(demux_data_in_62));
    InMux I__1295 (
            .O(N__11476),
            .I(N__11473));
    LocalMux I__1294 (
            .O(N__11473),
            .I(\demux.N_418_i_0_o2Z0Z_6 ));
    InMux I__1293 (
            .O(N__11470),
            .I(N__11467));
    LocalMux I__1292 (
            .O(N__11467),
            .I(N__11464));
    Span4Mux_h I__1291 (
            .O(N__11464),
            .I(N__11461));
    Span4Mux_h I__1290 (
            .O(N__11461),
            .I(N__11458));
    Span4Mux_v I__1289 (
            .O(N__11458),
            .I(N__11455));
    Odrv4 I__1288 (
            .O(N__11455),
            .I(demux_data_in_83));
    InMux I__1287 (
            .O(N__11452),
            .I(N__11449));
    LocalMux I__1286 (
            .O(N__11449),
            .I(demux_data_in_51));
    CascadeMux I__1285 (
            .O(N__11446),
            .I(\demux.N_835_cascade_ ));
    InMux I__1284 (
            .O(N__11443),
            .I(N__11440));
    LocalMux I__1283 (
            .O(N__11440),
            .I(demux_data_in_59));
    CascadeMux I__1282 (
            .O(N__11437),
            .I(N__11434));
    InMux I__1281 (
            .O(N__11434),
            .I(N__11431));
    LocalMux I__1280 (
            .O(N__11431),
            .I(N__11428));
    Odrv4 I__1279 (
            .O(N__11428),
            .I(demux_data_in_67));
    InMux I__1278 (
            .O(N__11425),
            .I(N__11422));
    LocalMux I__1277 (
            .O(N__11422),
            .I(\demux.N_421_i_0_o2Z0Z_6 ));
    InMux I__1276 (
            .O(N__11419),
            .I(N__11416));
    LocalMux I__1275 (
            .O(N__11416),
            .I(demux_data_in_63));
    InMux I__1274 (
            .O(N__11413),
            .I(N__11410));
    LocalMux I__1273 (
            .O(N__11410),
            .I(demux_data_in_57));
    InMux I__1272 (
            .O(N__11407),
            .I(N__11404));
    LocalMux I__1271 (
            .O(N__11404),
            .I(N__11401));
    Span4Mux_v I__1270 (
            .O(N__11401),
            .I(N__11398));
    Span4Mux_v I__1269 (
            .O(N__11398),
            .I(N__11395));
    Span4Mux_h I__1268 (
            .O(N__11395),
            .I(N__11392));
    Odrv4 I__1267 (
            .O(N__11392),
            .I(demux_data_in_87));
    InMux I__1266 (
            .O(N__11389),
            .I(N__11386));
    LocalMux I__1265 (
            .O(N__11386),
            .I(N__11383));
    Span4Mux_h I__1264 (
            .O(N__11383),
            .I(N__11380));
    Odrv4 I__1263 (
            .O(N__11380),
            .I(demux_data_in_79));
    CascadeMux I__1262 (
            .O(N__11377),
            .I(N__11373));
    CascadeMux I__1261 (
            .O(N__11376),
            .I(N__11370));
    InMux I__1260 (
            .O(N__11373),
            .I(N__11362));
    InMux I__1259 (
            .O(N__11370),
            .I(N__11362));
    InMux I__1258 (
            .O(N__11369),
            .I(N__11362));
    LocalMux I__1257 (
            .O(N__11362),
            .I(N__11359));
    Odrv4 I__1256 (
            .O(N__11359),
            .I(\sb_translator_1.N_1092 ));
    CascadeMux I__1255 (
            .O(N__11356),
            .I(\sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_ ));
    CEMux I__1254 (
            .O(N__11353),
            .I(N__11350));
    LocalMux I__1253 (
            .O(N__11350),
            .I(N__11347));
    Span4Mux_h I__1252 (
            .O(N__11347),
            .I(N__11344));
    Span4Mux_h I__1251 (
            .O(N__11344),
            .I(N__11341));
    Odrv4 I__1250 (
            .O(N__11341),
            .I(ram_we_11));
    CascadeMux I__1249 (
            .O(N__11338),
            .I(\sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_ ));
    InMux I__1248 (
            .O(N__11335),
            .I(N__11332));
    LocalMux I__1247 (
            .O(N__11332),
            .I(N__11325));
    InMux I__1246 (
            .O(N__11331),
            .I(N__11316));
    InMux I__1245 (
            .O(N__11330),
            .I(N__11316));
    InMux I__1244 (
            .O(N__11329),
            .I(N__11316));
    InMux I__1243 (
            .O(N__11328),
            .I(N__11316));
    Span4Mux_v I__1242 (
            .O(N__11325),
            .I(N__11313));
    LocalMux I__1241 (
            .O(N__11316),
            .I(N__11310));
    Span4Mux_v I__1240 (
            .O(N__11313),
            .I(N__11307));
    Span4Mux_v I__1239 (
            .O(N__11310),
            .I(N__11304));
    Odrv4 I__1238 (
            .O(N__11307),
            .I(mosi_data_out_17));
    Odrv4 I__1237 (
            .O(N__11304),
            .I(mosi_data_out_17));
    InMux I__1236 (
            .O(N__11299),
            .I(N__11296));
    LocalMux I__1235 (
            .O(N__11296),
            .I(N__11293));
    Span4Mux_v I__1234 (
            .O(N__11293),
            .I(N__11290));
    Span4Mux_v I__1233 (
            .O(N__11290),
            .I(N__11287));
    Span4Mux_h I__1232 (
            .O(N__11287),
            .I(N__11284));
    Odrv4 I__1231 (
            .O(N__11284),
            .I(demux_data_in_86));
    InMux I__1230 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__1229 (
            .O(N__11278),
            .I(N__11275));
    Span4Mux_v I__1228 (
            .O(N__11275),
            .I(N__11271));
    InMux I__1227 (
            .O(N__11274),
            .I(N__11268));
    Span4Mux_v I__1226 (
            .O(N__11271),
            .I(N__11265));
    LocalMux I__1225 (
            .O(N__11268),
            .I(N__11262));
    Span4Mux_h I__1224 (
            .O(N__11265),
            .I(N__11259));
    Span4Mux_h I__1223 (
            .O(N__11262),
            .I(N__11256));
    Span4Mux_h I__1222 (
            .O(N__11259),
            .I(N__11253));
    Span4Mux_h I__1221 (
            .O(N__11256),
            .I(N__11250));
    Odrv4 I__1220 (
            .O(N__11253),
            .I(reset_n));
    Odrv4 I__1219 (
            .O(N__11250),
            .I(reset_n));
    IoInMux I__1218 (
            .O(N__11245),
            .I(N__11242));
    LocalMux I__1217 (
            .O(N__11242),
            .I(N__11239));
    IoSpan4Mux I__1216 (
            .O(N__11239),
            .I(N__11236));
    Span4Mux_s3_v I__1215 (
            .O(N__11236),
            .I(N__11233));
    Odrv4 I__1214 (
            .O(N__11233),
            .I(reset_n_i));
    CEMux I__1213 (
            .O(N__11230),
            .I(N__11227));
    LocalMux I__1212 (
            .O(N__11227),
            .I(N__11224));
    Span4Mux_s2_v I__1211 (
            .O(N__11224),
            .I(N__11221));
    Span4Mux_h I__1210 (
            .O(N__11221),
            .I(N__11218));
    Odrv4 I__1209 (
            .O(N__11218),
            .I(ram_we_3));
    CEMux I__1208 (
            .O(N__11215),
            .I(N__11212));
    LocalMux I__1207 (
            .O(N__11212),
            .I(N__11209));
    Sp12to4 I__1206 (
            .O(N__11209),
            .I(N__11206));
    Span12Mux_s7_v I__1205 (
            .O(N__11206),
            .I(N__11203));
    Odrv12 I__1204 (
            .O(N__11203),
            .I(ram_we_13));
    CascadeMux I__1203 (
            .O(N__11200),
            .I(\sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_ ));
    CEMux I__1202 (
            .O(N__11197),
            .I(N__11194));
    LocalMux I__1201 (
            .O(N__11194),
            .I(ram_we_5));
    CEMux I__1200 (
            .O(N__11191),
            .I(N__11188));
    LocalMux I__1199 (
            .O(N__11188),
            .I(N__11185));
    Span4Mux_h I__1198 (
            .O(N__11185),
            .I(N__11182));
    Span4Mux_s0_h I__1197 (
            .O(N__11182),
            .I(N__11179));
    Span4Mux_h I__1196 (
            .O(N__11179),
            .I(N__11176));
    Odrv4 I__1195 (
            .O(N__11176),
            .I(ram_we_7));
    CEMux I__1194 (
            .O(N__11173),
            .I(N__11170));
    LocalMux I__1193 (
            .O(N__11170),
            .I(N__11167));
    Span12Mux_s7_v I__1192 (
            .O(N__11167),
            .I(N__11164));
    Odrv12 I__1191 (
            .O(N__11164),
            .I(ram_we_9));
    InMux I__1190 (
            .O(N__11161),
            .I(N__11158));
    LocalMux I__1189 (
            .O(N__11158),
            .I(N__11155));
    Span4Mux_v I__1188 (
            .O(N__11155),
            .I(N__11151));
    InMux I__1187 (
            .O(N__11154),
            .I(N__11148));
    Odrv4 I__1186 (
            .O(N__11151),
            .I(\spi_slave_1.mosi_data_inZ0Z_1 ));
    LocalMux I__1185 (
            .O(N__11148),
            .I(\spi_slave_1.mosi_data_inZ0Z_1 ));
    InMux I__1184 (
            .O(N__11143),
            .I(N__11140));
    LocalMux I__1183 (
            .O(N__11140),
            .I(N__11137));
    Odrv12 I__1182 (
            .O(N__11137),
            .I(\sb_translator_1.un1_num_leds_n_9 ));
    InMux I__1181 (
            .O(N__11134),
            .I(bfn_4_4_0_));
    InMux I__1180 (
            .O(N__11131),
            .I(N__11128));
    LocalMux I__1179 (
            .O(N__11128),
            .I(N__11125));
    Odrv12 I__1178 (
            .O(N__11125),
            .I(\sb_translator_1.un1_num_leds_n_10 ));
    InMux I__1177 (
            .O(N__11122),
            .I(\sb_translator_1.un1_num_leds_0_cry_9 ));
    CascadeMux I__1176 (
            .O(N__11119),
            .I(N__11116));
    InMux I__1175 (
            .O(N__11116),
            .I(N__11113));
    LocalMux I__1174 (
            .O(N__11113),
            .I(N__11110));
    Odrv4 I__1173 (
            .O(N__11110),
            .I(\sb_translator_1.un1_num_leds_n_11 ));
    InMux I__1172 (
            .O(N__11107),
            .I(\sb_translator_1.un1_num_leds_0_cry_10 ));
    InMux I__1171 (
            .O(N__11104),
            .I(N__11101));
    LocalMux I__1170 (
            .O(N__11101),
            .I(N__11098));
    Odrv4 I__1169 (
            .O(N__11098),
            .I(\sb_translator_1.un1_num_leds_n_12 ));
    InMux I__1168 (
            .O(N__11095),
            .I(\sb_translator_1.un1_num_leds_0_cry_11 ));
    InMux I__1167 (
            .O(N__11092),
            .I(N__11089));
    LocalMux I__1166 (
            .O(N__11089),
            .I(N__11086));
    Odrv4 I__1165 (
            .O(N__11086),
            .I(\sb_translator_1.un1_num_leds_n_13 ));
    InMux I__1164 (
            .O(N__11083),
            .I(\sb_translator_1.un1_num_leds_0_cry_12 ));
    InMux I__1163 (
            .O(N__11080),
            .I(N__11077));
    LocalMux I__1162 (
            .O(N__11077),
            .I(N__11074));
    Odrv4 I__1161 (
            .O(N__11074),
            .I(\sb_translator_1.un1_num_leds_n_14 ));
    InMux I__1160 (
            .O(N__11071),
            .I(\sb_translator_1.un1_num_leds_0_cry_13 ));
    InMux I__1159 (
            .O(N__11068),
            .I(N__11065));
    LocalMux I__1158 (
            .O(N__11065),
            .I(N__11062));
    Odrv4 I__1157 (
            .O(N__11062),
            .I(\sb_translator_1.un1_num_leds_n_15 ));
    InMux I__1156 (
            .O(N__11059),
            .I(\sb_translator_1.un1_num_leds_0_cry_14 ));
    InMux I__1155 (
            .O(N__11056),
            .I(\sb_translator_1.un1_num_leds_0_cry_15 ));
    InMux I__1154 (
            .O(N__11053),
            .I(N__11050));
    LocalMux I__1153 (
            .O(N__11050),
            .I(N__11047));
    Span4Mux_h I__1152 (
            .O(N__11047),
            .I(N__11044));
    Odrv4 I__1151 (
            .O(N__11044),
            .I(\sb_translator_1.un1_num_leds_n_16 ));
    InMux I__1150 (
            .O(N__11041),
            .I(N__11038));
    LocalMux I__1149 (
            .O(N__11038),
            .I(N__11035));
    Odrv12 I__1148 (
            .O(N__11035),
            .I(\sb_translator_1.un1_num_leds_n_1 ));
    InMux I__1147 (
            .O(N__11032),
            .I(N__11029));
    LocalMux I__1146 (
            .O(N__11029),
            .I(N__11026));
    Odrv12 I__1145 (
            .O(N__11026),
            .I(\sb_translator_1.un1_num_leds_n_2 ));
    InMux I__1144 (
            .O(N__11023),
            .I(\sb_translator_1.un1_num_leds_0_cry_1 ));
    CascadeMux I__1143 (
            .O(N__11020),
            .I(N__11017));
    InMux I__1142 (
            .O(N__11017),
            .I(N__11014));
    LocalMux I__1141 (
            .O(N__11014),
            .I(N__11011));
    Odrv4 I__1140 (
            .O(N__11011),
            .I(\sb_translator_1.un1_num_leds_n_3 ));
    InMux I__1139 (
            .O(N__11008),
            .I(\sb_translator_1.un1_num_leds_0_cry_2 ));
    InMux I__1138 (
            .O(N__11005),
            .I(N__11002));
    LocalMux I__1137 (
            .O(N__11002),
            .I(N__10999));
    Odrv4 I__1136 (
            .O(N__10999),
            .I(\sb_translator_1.un1_num_leds_n_4 ));
    InMux I__1135 (
            .O(N__10996),
            .I(\sb_translator_1.un1_num_leds_0_cry_3 ));
    InMux I__1134 (
            .O(N__10993),
            .I(N__10990));
    LocalMux I__1133 (
            .O(N__10990),
            .I(N__10987));
    Odrv4 I__1132 (
            .O(N__10987),
            .I(\sb_translator_1.un1_num_leds_n_5 ));
    InMux I__1131 (
            .O(N__10984),
            .I(\sb_translator_1.un1_num_leds_0_cry_4 ));
    CascadeMux I__1130 (
            .O(N__10981),
            .I(N__10978));
    InMux I__1129 (
            .O(N__10978),
            .I(N__10975));
    LocalMux I__1128 (
            .O(N__10975),
            .I(N__10972));
    Odrv4 I__1127 (
            .O(N__10972),
            .I(\sb_translator_1.un1_num_leds_n_6 ));
    InMux I__1126 (
            .O(N__10969),
            .I(\sb_translator_1.un1_num_leds_0_cry_5 ));
    InMux I__1125 (
            .O(N__10966),
            .I(N__10963));
    LocalMux I__1124 (
            .O(N__10963),
            .I(N__10960));
    Odrv4 I__1123 (
            .O(N__10960),
            .I(\sb_translator_1.un1_num_leds_n_7 ));
    InMux I__1122 (
            .O(N__10957),
            .I(\sb_translator_1.un1_num_leds_0_cry_6 ));
    InMux I__1121 (
            .O(N__10954),
            .I(N__10951));
    LocalMux I__1120 (
            .O(N__10951),
            .I(N__10948));
    Span4Mux_h I__1119 (
            .O(N__10948),
            .I(N__10945));
    Odrv4 I__1118 (
            .O(N__10945),
            .I(\sb_translator_1.un1_num_leds_n_8 ));
    InMux I__1117 (
            .O(N__10942),
            .I(\sb_translator_1.un1_num_leds_0_cry_7 ));
    CascadeMux I__1116 (
            .O(N__10939),
            .I(\spi_slave_1.N_49_0_cascade_ ));
    CascadeMux I__1115 (
            .O(N__10936),
            .I(\spi_slave_1.N_25_0_cascade_ ));
    InMux I__1114 (
            .O(N__10933),
            .I(N__10930));
    LocalMux I__1113 (
            .O(N__10930),
            .I(N__10927));
    Span4Mux_s3_h I__1112 (
            .O(N__10927),
            .I(N__10924));
    Odrv4 I__1111 (
            .O(N__10924),
            .I(\spi_slave_1.miso_data_outZ0Z_23 ));
    CascadeMux I__1110 (
            .O(N__10921),
            .I(N__10916));
    InMux I__1109 (
            .O(N__10920),
            .I(N__10911));
    InMux I__1108 (
            .O(N__10919),
            .I(N__10908));
    InMux I__1107 (
            .O(N__10916),
            .I(N__10901));
    InMux I__1106 (
            .O(N__10915),
            .I(N__10901));
    InMux I__1105 (
            .O(N__10914),
            .I(N__10901));
    LocalMux I__1104 (
            .O(N__10911),
            .I(N__10898));
    LocalMux I__1103 (
            .O(N__10908),
            .I(\spi_slave_1.miso_data_out_0_sqmuxa ));
    LocalMux I__1102 (
            .O(N__10901),
            .I(\spi_slave_1.miso_data_out_0_sqmuxa ));
    Odrv4 I__1101 (
            .O(N__10898),
            .I(\spi_slave_1.miso_data_out_0_sqmuxa ));
    InMux I__1100 (
            .O(N__10891),
            .I(N__10888));
    LocalMux I__1099 (
            .O(N__10888),
            .I(\spi_slave_1.N_96_mux ));
    InMux I__1098 (
            .O(N__10885),
            .I(N__10880));
    InMux I__1097 (
            .O(N__10884),
            .I(N__10877));
    InMux I__1096 (
            .O(N__10883),
            .I(N__10874));
    LocalMux I__1095 (
            .O(N__10880),
            .I(\spi_slave_1.N_94_mux ));
    LocalMux I__1094 (
            .O(N__10877),
            .I(\spi_slave_1.N_94_mux ));
    LocalMux I__1093 (
            .O(N__10874),
            .I(\spi_slave_1.N_94_mux ));
    CascadeMux I__1092 (
            .O(N__10867),
            .I(\spi_slave_1.N_94_mux_cascade_ ));
    InMux I__1091 (
            .O(N__10864),
            .I(N__10852));
    InMux I__1090 (
            .O(N__10863),
            .I(N__10852));
    InMux I__1089 (
            .O(N__10862),
            .I(N__10852));
    InMux I__1088 (
            .O(N__10861),
            .I(N__10849));
    InMux I__1087 (
            .O(N__10860),
            .I(N__10846));
    InMux I__1086 (
            .O(N__10859),
            .I(N__10843));
    LocalMux I__1085 (
            .O(N__10852),
            .I(N__10840));
    LocalMux I__1084 (
            .O(N__10849),
            .I(\spi_slave_1.bitcnt_txZ0Z_3 ));
    LocalMux I__1083 (
            .O(N__10846),
            .I(\spi_slave_1.bitcnt_txZ0Z_3 ));
    LocalMux I__1082 (
            .O(N__10843),
            .I(\spi_slave_1.bitcnt_txZ0Z_3 ));
    Odrv4 I__1081 (
            .O(N__10840),
            .I(\spi_slave_1.bitcnt_txZ0Z_3 ));
    InMux I__1080 (
            .O(N__10831),
            .I(N__10825));
    InMux I__1079 (
            .O(N__10830),
            .I(N__10825));
    LocalMux I__1078 (
            .O(N__10825),
            .I(\spi_slave_1.N_17_0 ));
    InMux I__1077 (
            .O(N__10822),
            .I(N__10819));
    LocalMux I__1076 (
            .O(N__10819),
            .I(\spi_slave_1.N_20_0 ));
    InMux I__1075 (
            .O(N__10816),
            .I(N__10813));
    LocalMux I__1074 (
            .O(N__10813),
            .I(\spi_slave_1.N_91 ));
    IoInMux I__1073 (
            .O(N__10810),
            .I(N__10807));
    LocalMux I__1072 (
            .O(N__10807),
            .I(N__10803));
    InMux I__1071 (
            .O(N__10806),
            .I(N__10800));
    Odrv4 I__1070 (
            .O(N__10803),
            .I(miso));
    LocalMux I__1069 (
            .O(N__10800),
            .I(miso));
    IoInMux I__1068 (
            .O(N__10795),
            .I(N__10792));
    LocalMux I__1067 (
            .O(N__10792),
            .I(N__10789));
    IoSpan4Mux I__1066 (
            .O(N__10789),
            .I(N__10786));
    Odrv4 I__1065 (
            .O(N__10786),
            .I(\spi_slave_1.bitcnt_rxe_0_i ));
    CascadeMux I__1064 (
            .O(N__10783),
            .I(N__10780));
    InMux I__1063 (
            .O(N__10780),
            .I(N__10777));
    LocalMux I__1062 (
            .O(N__10777),
            .I(\spi_slave_1.bitcnt_tx10 ));
    CascadeMux I__1061 (
            .O(N__10774),
            .I(\spi_slave_1.bitcnt_tx10_cascade_ ));
    InMux I__1060 (
            .O(N__10771),
            .I(N__10768));
    LocalMux I__1059 (
            .O(N__10768),
            .I(N__10765));
    Odrv4 I__1058 (
            .O(N__10765),
            .I(\spi_slave_1.miso_data_outZ0Z_8 ));
    InMux I__1057 (
            .O(N__10762),
            .I(N__10758));
    InMux I__1056 (
            .O(N__10761),
            .I(N__10755));
    LocalMux I__1055 (
            .O(N__10758),
            .I(N__10752));
    LocalMux I__1054 (
            .O(N__10755),
            .I(N__10747));
    Span4Mux_v I__1053 (
            .O(N__10752),
            .I(N__10747));
    Odrv4 I__1052 (
            .O(N__10747),
            .I(miso_tx));
    InMux I__1051 (
            .O(N__10744),
            .I(N__10741));
    LocalMux I__1050 (
            .O(N__10741),
            .I(N__10738));
    Odrv4 I__1049 (
            .O(N__10738),
            .I(\spi_slave_1.N_82 ));
    InMux I__1048 (
            .O(N__10735),
            .I(N__10732));
    LocalMux I__1047 (
            .O(N__10732),
            .I(\spi_slave_1.miso_RNOZ0Z_17 ));
    InMux I__1046 (
            .O(N__10729),
            .I(N__10726));
    LocalMux I__1045 (
            .O(N__10726),
            .I(N__10723));
    Odrv4 I__1044 (
            .O(N__10723),
            .I(\spi_slave_1.miso_RNOZ0Z_10 ));
    CascadeMux I__1043 (
            .O(N__10720),
            .I(\spi_slave_1.m48_ns_1_cascade_ ));
    InMux I__1042 (
            .O(N__10717),
            .I(N__10714));
    LocalMux I__1041 (
            .O(N__10714),
            .I(miso_data_in_8));
    InMux I__1040 (
            .O(N__10711),
            .I(N__10705));
    InMux I__1039 (
            .O(N__10710),
            .I(N__10705));
    LocalMux I__1038 (
            .O(N__10705),
            .I(N__10699));
    InMux I__1037 (
            .O(N__10704),
            .I(N__10692));
    InMux I__1036 (
            .O(N__10703),
            .I(N__10692));
    InMux I__1035 (
            .O(N__10702),
            .I(N__10692));
    Odrv4 I__1034 (
            .O(N__10699),
            .I(\spi_slave_1.clk_pos_i ));
    LocalMux I__1033 (
            .O(N__10692),
            .I(\spi_slave_1.clk_pos_i ));
    CascadeMux I__1032 (
            .O(N__10687),
            .I(N__10684));
    InMux I__1031 (
            .O(N__10684),
            .I(N__10681));
    LocalMux I__1030 (
            .O(N__10681),
            .I(\spi_slave_1.miso_data_outZ0Z_22 ));
    InMux I__1029 (
            .O(N__10678),
            .I(N__10675));
    LocalMux I__1028 (
            .O(N__10675),
            .I(\spi_slave_1.miso_data_outZ0Z_21 ));
    CascadeMux I__1027 (
            .O(N__10672),
            .I(\spi_slave_1.m81_ns_1_cascade_ ));
    InMux I__1026 (
            .O(N__10669),
            .I(N__10666));
    LocalMux I__1025 (
            .O(N__10666),
            .I(\spi_slave_1.miso_data_outZ0Z_5 ));
    InMux I__1024 (
            .O(N__10663),
            .I(N__10660));
    LocalMux I__1023 (
            .O(N__10660),
            .I(\spi_slave_1.miso_data_outZ0Z_4 ));
    CascadeMux I__1022 (
            .O(N__10657),
            .I(N__10654));
    InMux I__1021 (
            .O(N__10654),
            .I(N__10651));
    LocalMux I__1020 (
            .O(N__10651),
            .I(\spi_slave_1.miso_data_outZ0Z_20 ));
    InMux I__1019 (
            .O(N__10648),
            .I(N__10645));
    LocalMux I__1018 (
            .O(N__10645),
            .I(\spi_slave_1.miso_data_outZ0Z_19 ));
    CascadeMux I__1017 (
            .O(N__10642),
            .I(\spi_slave_1.m60_ns_1_cascade_ ));
    InMux I__1016 (
            .O(N__10639),
            .I(N__10636));
    LocalMux I__1015 (
            .O(N__10636),
            .I(N__10633));
    Odrv12 I__1014 (
            .O(N__10633),
            .I(clk_spi));
    CascadeMux I__1013 (
            .O(N__10630),
            .I(N__10626));
    InMux I__1012 (
            .O(N__10629),
            .I(N__10623));
    InMux I__1011 (
            .O(N__10626),
            .I(N__10620));
    LocalMux I__1010 (
            .O(N__10623),
            .I(\sb_translator_1.instr_tmpZ0Z_22 ));
    LocalMux I__1009 (
            .O(N__10620),
            .I(\sb_translator_1.instr_tmpZ0Z_22 ));
    CascadeMux I__1008 (
            .O(N__10615),
            .I(N__10611));
    InMux I__1007 (
            .O(N__10614),
            .I(N__10608));
    InMux I__1006 (
            .O(N__10611),
            .I(N__10605));
    LocalMux I__1005 (
            .O(N__10608),
            .I(\sb_translator_1.instr_tmpZ0Z_23 ));
    LocalMux I__1004 (
            .O(N__10605),
            .I(\sb_translator_1.instr_tmpZ0Z_23 ));
    InMux I__1003 (
            .O(N__10600),
            .I(N__10597));
    LocalMux I__1002 (
            .O(N__10597),
            .I(miso_data_in_19));
    InMux I__1001 (
            .O(N__10594),
            .I(N__10591));
    LocalMux I__1000 (
            .O(N__10591),
            .I(miso_data_in_20));
    InMux I__999 (
            .O(N__10588),
            .I(N__10585));
    LocalMux I__998 (
            .O(N__10585),
            .I(miso_data_in_21));
    InMux I__997 (
            .O(N__10582),
            .I(N__10579));
    LocalMux I__996 (
            .O(N__10579),
            .I(miso_data_in_22));
    InMux I__995 (
            .O(N__10576),
            .I(N__10573));
    LocalMux I__994 (
            .O(N__10573),
            .I(miso_data_in_23));
    InMux I__993 (
            .O(N__10570),
            .I(N__10567));
    LocalMux I__992 (
            .O(N__10567),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_9 ));
    InMux I__991 (
            .O(N__10564),
            .I(N__10561));
    LocalMux I__990 (
            .O(N__10561),
            .I(N__10553));
    InMux I__989 (
            .O(N__10560),
            .I(N__10544));
    InMux I__988 (
            .O(N__10559),
            .I(N__10544));
    InMux I__987 (
            .O(N__10558),
            .I(N__10544));
    InMux I__986 (
            .O(N__10557),
            .I(N__10544));
    InMux I__985 (
            .O(N__10556),
            .I(N__10541));
    Span4Mux_s2_h I__984 (
            .O(N__10553),
            .I(N__10538));
    LocalMux I__983 (
            .O(N__10544),
            .I(\sb_translator_1.cntZ0Z_9 ));
    LocalMux I__982 (
            .O(N__10541),
            .I(\sb_translator_1.cntZ0Z_9 ));
    Odrv4 I__981 (
            .O(N__10538),
            .I(\sb_translator_1.cntZ0Z_9 ));
    InMux I__980 (
            .O(N__10531),
            .I(N__10526));
    CascadeMux I__979 (
            .O(N__10530),
            .I(N__10523));
    CascadeMux I__978 (
            .O(N__10529),
            .I(N__10519));
    LocalMux I__977 (
            .O(N__10526),
            .I(N__10514));
    InMux I__976 (
            .O(N__10523),
            .I(N__10505));
    InMux I__975 (
            .O(N__10522),
            .I(N__10505));
    InMux I__974 (
            .O(N__10519),
            .I(N__10505));
    InMux I__973 (
            .O(N__10518),
            .I(N__10505));
    InMux I__972 (
            .O(N__10517),
            .I(N__10502));
    Span4Mux_s2_h I__971 (
            .O(N__10514),
            .I(N__10499));
    LocalMux I__970 (
            .O(N__10505),
            .I(\sb_translator_1.cntZ0Z_12 ));
    LocalMux I__969 (
            .O(N__10502),
            .I(\sb_translator_1.cntZ0Z_12 ));
    Odrv4 I__968 (
            .O(N__10499),
            .I(\sb_translator_1.cntZ0Z_12 ));
    CascadeMux I__967 (
            .O(N__10492),
            .I(N__10488));
    InMux I__966 (
            .O(N__10491),
            .I(N__10485));
    InMux I__965 (
            .O(N__10488),
            .I(N__10482));
    LocalMux I__964 (
            .O(N__10485),
            .I(\sb_translator_1.instr_tmpZ0Z_18 ));
    LocalMux I__963 (
            .O(N__10482),
            .I(\sb_translator_1.instr_tmpZ0Z_18 ));
    CascadeMux I__962 (
            .O(N__10477),
            .I(N__10473));
    InMux I__961 (
            .O(N__10476),
            .I(N__10470));
    InMux I__960 (
            .O(N__10473),
            .I(N__10467));
    LocalMux I__959 (
            .O(N__10470),
            .I(\sb_translator_1.instr_tmpZ0Z_19 ));
    LocalMux I__958 (
            .O(N__10467),
            .I(\sb_translator_1.instr_tmpZ0Z_19 ));
    CascadeMux I__957 (
            .O(N__10462),
            .I(N__10458));
    InMux I__956 (
            .O(N__10461),
            .I(N__10455));
    InMux I__955 (
            .O(N__10458),
            .I(N__10452));
    LocalMux I__954 (
            .O(N__10455),
            .I(\sb_translator_1.instr_tmpZ0Z_20 ));
    LocalMux I__953 (
            .O(N__10452),
            .I(\sb_translator_1.instr_tmpZ0Z_20 ));
    CascadeMux I__952 (
            .O(N__10447),
            .I(N__10443));
    InMux I__951 (
            .O(N__10446),
            .I(N__10440));
    InMux I__950 (
            .O(N__10443),
            .I(N__10437));
    LocalMux I__949 (
            .O(N__10440),
            .I(\sb_translator_1.instr_tmpZ0Z_21 ));
    LocalMux I__948 (
            .O(N__10437),
            .I(\sb_translator_1.instr_tmpZ0Z_21 ));
    CascadeMux I__947 (
            .O(N__10432),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_0_cascade_ ));
    InMux I__946 (
            .O(N__10429),
            .I(N__10426));
    LocalMux I__945 (
            .O(N__10426),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_13 ));
    InMux I__944 (
            .O(N__10423),
            .I(N__10419));
    InMux I__943 (
            .O(N__10422),
            .I(N__10416));
    LocalMux I__942 (
            .O(N__10419),
            .I(N__10413));
    LocalMux I__941 (
            .O(N__10416),
            .I(\sb_translator_1.cntZ0Z_13 ));
    Odrv4 I__940 (
            .O(N__10413),
            .I(\sb_translator_1.cntZ0Z_13 ));
    InMux I__939 (
            .O(N__10408),
            .I(N__10405));
    LocalMux I__938 (
            .O(N__10405),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_14 ));
    InMux I__937 (
            .O(N__10402),
            .I(N__10398));
    InMux I__936 (
            .O(N__10401),
            .I(N__10395));
    LocalMux I__935 (
            .O(N__10398),
            .I(N__10392));
    LocalMux I__934 (
            .O(N__10395),
            .I(\sb_translator_1.cntZ0Z_14 ));
    Odrv4 I__933 (
            .O(N__10392),
            .I(\sb_translator_1.cntZ0Z_14 ));
    InMux I__932 (
            .O(N__10387),
            .I(N__10384));
    LocalMux I__931 (
            .O(N__10384),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_15 ));
    InMux I__930 (
            .O(N__10381),
            .I(N__10377));
    InMux I__929 (
            .O(N__10380),
            .I(N__10374));
    LocalMux I__928 (
            .O(N__10377),
            .I(N__10371));
    LocalMux I__927 (
            .O(N__10374),
            .I(\sb_translator_1.cntZ0Z_15 ));
    Odrv4 I__926 (
            .O(N__10371),
            .I(\sb_translator_1.cntZ0Z_15 ));
    InMux I__925 (
            .O(N__10366),
            .I(N__10363));
    LocalMux I__924 (
            .O(N__10363),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_16 ));
    InMux I__923 (
            .O(N__10360),
            .I(N__10356));
    InMux I__922 (
            .O(N__10359),
            .I(N__10353));
    LocalMux I__921 (
            .O(N__10356),
            .I(\sb_translator_1.cntZ0Z_16 ));
    LocalMux I__920 (
            .O(N__10353),
            .I(\sb_translator_1.cntZ0Z_16 ));
    InMux I__919 (
            .O(N__10348),
            .I(N__10345));
    LocalMux I__918 (
            .O(N__10345),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_1 ));
    InMux I__917 (
            .O(N__10342),
            .I(N__10339));
    LocalMux I__916 (
            .O(N__10339),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_11 ));
    InMux I__915 (
            .O(N__10336),
            .I(N__10333));
    LocalMux I__914 (
            .O(N__10333),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_12 ));
    InMux I__913 (
            .O(N__10330),
            .I(N__10327));
    LocalMux I__912 (
            .O(N__10327),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_10 ));
    InMux I__911 (
            .O(N__10324),
            .I(N__10321));
    LocalMux I__910 (
            .O(N__10321),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_2 ));
    InMux I__909 (
            .O(N__10318),
            .I(N__10315));
    LocalMux I__908 (
            .O(N__10315),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_3 ));
    InMux I__907 (
            .O(N__10312),
            .I(N__10309));
    LocalMux I__906 (
            .O(N__10309),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_4 ));
    InMux I__905 (
            .O(N__10306),
            .I(N__10303));
    LocalMux I__904 (
            .O(N__10303),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_5 ));
    InMux I__903 (
            .O(N__10300),
            .I(N__10297));
    LocalMux I__902 (
            .O(N__10297),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_6 ));
    InMux I__901 (
            .O(N__10294),
            .I(N__10291));
    LocalMux I__900 (
            .O(N__10291),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_7 ));
    InMux I__899 (
            .O(N__10288),
            .I(N__10285));
    LocalMux I__898 (
            .O(N__10285),
            .I(\sb_translator_1.cnt_RNO_0Z0Z_8 ));
    InMux I__897 (
            .O(N__10282),
            .I(N__10278));
    InMux I__896 (
            .O(N__10281),
            .I(N__10275));
    LocalMux I__895 (
            .O(N__10278),
            .I(\sb_translator_1.stateZ0Z_5 ));
    LocalMux I__894 (
            .O(N__10275),
            .I(\sb_translator_1.stateZ0Z_5 ));
    InMux I__893 (
            .O(N__10270),
            .I(N__10267));
    LocalMux I__892 (
            .O(N__10267),
            .I(\spi_slave_1.mosi_data_inZ0Z_23 ));
    InMux I__891 (
            .O(N__10264),
            .I(N__10260));
    InMux I__890 (
            .O(N__10263),
            .I(N__10257));
    LocalMux I__889 (
            .O(N__10260),
            .I(\spi_slave_1.mosi_data_inZ0Z_18 ));
    LocalMux I__888 (
            .O(N__10257),
            .I(\spi_slave_1.mosi_data_inZ0Z_18 ));
    InMux I__887 (
            .O(N__10252),
            .I(N__10248));
    InMux I__886 (
            .O(N__10251),
            .I(N__10245));
    LocalMux I__885 (
            .O(N__10248),
            .I(\spi_slave_1.mosi_data_inZ0Z_19 ));
    LocalMux I__884 (
            .O(N__10245),
            .I(\spi_slave_1.mosi_data_inZ0Z_19 ));
    InMux I__883 (
            .O(N__10240),
            .I(N__10236));
    InMux I__882 (
            .O(N__10239),
            .I(N__10233));
    LocalMux I__881 (
            .O(N__10236),
            .I(\spi_slave_1.mosi_data_inZ0Z_20 ));
    LocalMux I__880 (
            .O(N__10233),
            .I(\spi_slave_1.mosi_data_inZ0Z_20 ));
    InMux I__879 (
            .O(N__10228),
            .I(N__10224));
    InMux I__878 (
            .O(N__10227),
            .I(N__10221));
    LocalMux I__877 (
            .O(N__10224),
            .I(\spi_slave_1.mosi_data_inZ0Z_21 ));
    LocalMux I__876 (
            .O(N__10221),
            .I(\spi_slave_1.mosi_data_inZ0Z_21 ));
    InMux I__875 (
            .O(N__10216),
            .I(N__10212));
    InMux I__874 (
            .O(N__10215),
            .I(N__10209));
    LocalMux I__873 (
            .O(N__10212),
            .I(\spi_slave_1.mosi_data_inZ0Z_22 ));
    LocalMux I__872 (
            .O(N__10209),
            .I(\spi_slave_1.mosi_data_inZ0Z_22 ));
    InMux I__871 (
            .O(N__10204),
            .I(N__10201));
    LocalMux I__870 (
            .O(N__10201),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO ));
    InMux I__869 (
            .O(N__10198),
            .I(N__10195));
    LocalMux I__868 (
            .O(N__10195),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO ));
    InMux I__867 (
            .O(N__10192),
            .I(N__10188));
    InMux I__866 (
            .O(N__10191),
            .I(N__10185));
    LocalMux I__865 (
            .O(N__10188),
            .I(\spi_slave_1.bitcnt_rxZ0Z_3 ));
    LocalMux I__864 (
            .O(N__10185),
            .I(\spi_slave_1.bitcnt_rxZ0Z_3 ));
    InMux I__863 (
            .O(N__10180),
            .I(\spi_slave_1.bitcnt_rx_cry_2 ));
    InMux I__862 (
            .O(N__10177),
            .I(\spi_slave_1.bitcnt_rx_cry_3 ));
    InMux I__861 (
            .O(N__10174),
            .I(N__10169));
    InMux I__860 (
            .O(N__10173),
            .I(N__10164));
    InMux I__859 (
            .O(N__10172),
            .I(N__10164));
    LocalMux I__858 (
            .O(N__10169),
            .I(\spi_slave_1.bitcnt_rxZ0Z_4 ));
    LocalMux I__857 (
            .O(N__10164),
            .I(\spi_slave_1.bitcnt_rxZ0Z_4 ));
    InMux I__856 (
            .O(N__10159),
            .I(N__10156));
    LocalMux I__855 (
            .O(N__10156),
            .I(miso_en));
    InMux I__854 (
            .O(N__10153),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_0 ));
    InMux I__853 (
            .O(N__10150),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_1 ));
    InMux I__852 (
            .O(N__10147),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_2 ));
    InMux I__851 (
            .O(N__10144),
            .I(\spi_slave_1.un1_bitcnt_tx_1_cry_3 ));
    InMux I__850 (
            .O(N__10141),
            .I(N__10138));
    LocalMux I__849 (
            .O(N__10138),
            .I(\spi_slave_1.un3_mosi_data_out_3 ));
    CascadeMux I__848 (
            .O(N__10135),
            .I(\spi_slave_1.un3_mosi_data_out_3_cascade_ ));
    InMux I__847 (
            .O(N__10132),
            .I(N__10127));
    InMux I__846 (
            .O(N__10131),
            .I(N__10122));
    InMux I__845 (
            .O(N__10130),
            .I(N__10122));
    LocalMux I__844 (
            .O(N__10127),
            .I(\spi_slave_1.bitcnt_rxZ0Z_0 ));
    LocalMux I__843 (
            .O(N__10122),
            .I(\spi_slave_1.bitcnt_rxZ0Z_0 ));
    InMux I__842 (
            .O(N__10117),
            .I(bfn_1_10_0_));
    InMux I__841 (
            .O(N__10114),
            .I(N__10110));
    InMux I__840 (
            .O(N__10113),
            .I(N__10107));
    LocalMux I__839 (
            .O(N__10110),
            .I(\spi_slave_1.bitcnt_rxZ0Z_1 ));
    LocalMux I__838 (
            .O(N__10107),
            .I(\spi_slave_1.bitcnt_rxZ0Z_1 ));
    InMux I__837 (
            .O(N__10102),
            .I(\spi_slave_1.bitcnt_rx_cry_0 ));
    InMux I__836 (
            .O(N__10099),
            .I(N__10095));
    InMux I__835 (
            .O(N__10098),
            .I(N__10092));
    LocalMux I__834 (
            .O(N__10095),
            .I(\spi_slave_1.bitcnt_rxZ0Z_2 ));
    LocalMux I__833 (
            .O(N__10092),
            .I(\spi_slave_1.bitcnt_rxZ0Z_2 ));
    InMux I__832 (
            .O(N__10087),
            .I(\spi_slave_1.bitcnt_rx_cry_1 ));
    InMux I__831 (
            .O(N__10084),
            .I(\sb_translator_1.cnt19_cry_31 ));
    InMux I__830 (
            .O(N__10081),
            .I(\sb_translator_1.cnt19_cry_32 ));
    InMux I__829 (
            .O(N__10078),
            .I(bfn_1_7_0_));
    InMux I__828 (
            .O(N__10075),
            .I(\sb_translator_1.cnt19_cry_34 ));
    InMux I__827 (
            .O(N__10072),
            .I(\sb_translator_1.cnt19_cry_35 ));
    IoInMux I__826 (
            .O(N__10069),
            .I(N__10066));
    LocalMux I__825 (
            .O(N__10066),
            .I(N__10063));
    Span4Mux_s1_v I__824 (
            .O(N__10063),
            .I(N__10060));
    Span4Mux_v I__823 (
            .O(N__10060),
            .I(N__10057));
    Odrv4 I__822 (
            .O(N__10057),
            .I(\spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4 ));
    InMux I__821 (
            .O(N__10054),
            .I(\sb_translator_1.cnt19_cry_22 ));
    InMux I__820 (
            .O(N__10051),
            .I(\sb_translator_1.cnt19_cry_23 ));
    InMux I__819 (
            .O(N__10048),
            .I(\sb_translator_1.cnt19_cry_24 ));
    InMux I__818 (
            .O(N__10045),
            .I(bfn_1_6_0_));
    InMux I__817 (
            .O(N__10042),
            .I(\sb_translator_1.cnt19_cry_26 ));
    InMux I__816 (
            .O(N__10039),
            .I(\sb_translator_1.cnt19_cry_27 ));
    InMux I__815 (
            .O(N__10036),
            .I(\sb_translator_1.cnt19_cry_28 ));
    InMux I__814 (
            .O(N__10033),
            .I(\sb_translator_1.cnt19_cry_29 ));
    InMux I__813 (
            .O(N__10030),
            .I(\sb_translator_1.cnt19_cry_30 ));
    CascadeMux I__812 (
            .O(N__10027),
            .I(N__10024));
    InMux I__811 (
            .O(N__10024),
            .I(N__10021));
    LocalMux I__810 (
            .O(N__10021),
            .I(N__10018));
    Odrv4 I__809 (
            .O(N__10018),
            .I(\sb_translator_1.cnt_RNI0G0QZ0Z_13 ));
    CascadeMux I__808 (
            .O(N__10015),
            .I(N__10012));
    InMux I__807 (
            .O(N__10012),
            .I(N__10009));
    LocalMux I__806 (
            .O(N__10009),
            .I(N__10006));
    Odrv4 I__805 (
            .O(N__10006),
            .I(\sb_translator_1.cnt_RNI4L1QZ0Z_14 ));
    CascadeMux I__804 (
            .O(N__10003),
            .I(N__10000));
    InMux I__803 (
            .O(N__10000),
            .I(N__9997));
    LocalMux I__802 (
            .O(N__9997),
            .I(N__9994));
    Odrv4 I__801 (
            .O(N__9994),
            .I(\sb_translator_1.cnt_RNI8Q2QZ0Z_15 ));
    CascadeMux I__800 (
            .O(N__9991),
            .I(N__9988));
    InMux I__799 (
            .O(N__9988),
            .I(N__9985));
    LocalMux I__798 (
            .O(N__9985),
            .I(\sb_translator_1.cnt_i_16 ));
    InMux I__797 (
            .O(N__9982),
            .I(\sb_translator_1.cnt19_cry_16 ));
    InMux I__796 (
            .O(N__9979),
            .I(\sb_translator_1.cnt19_cry_18 ));
    InMux I__795 (
            .O(N__9976),
            .I(\sb_translator_1.cnt19_cry_20 ));
    InMux I__794 (
            .O(N__9973),
            .I(\sb_translator_1.cnt19_cry_21 ));
    CascadeMux I__793 (
            .O(N__9970),
            .I(N__9967));
    InMux I__792 (
            .O(N__9967),
            .I(N__9964));
    LocalMux I__791 (
            .O(N__9964),
            .I(\sb_translator_1.cnt_RNI0T5OZ0Z_4 ));
    CascadeMux I__790 (
            .O(N__9961),
            .I(N__9958));
    InMux I__789 (
            .O(N__9958),
            .I(N__9955));
    LocalMux I__788 (
            .O(N__9955),
            .I(\sb_translator_1.cnt_RNI427OZ0Z_5 ));
    InMux I__787 (
            .O(N__9952),
            .I(N__9949));
    LocalMux I__786 (
            .O(N__9949),
            .I(\sb_translator_1.cnt_RNI878OZ0Z_6 ));
    CascadeMux I__785 (
            .O(N__9946),
            .I(N__9943));
    InMux I__784 (
            .O(N__9943),
            .I(N__9940));
    LocalMux I__783 (
            .O(N__9940),
            .I(\sb_translator_1.cnt_RNICC9OZ0Z_7 ));
    CascadeMux I__782 (
            .O(N__9937),
            .I(N__9934));
    InMux I__781 (
            .O(N__9934),
            .I(N__9931));
    LocalMux I__780 (
            .O(N__9931),
            .I(\sb_translator_1.cnt_RNIGHAOZ0Z_8 ));
    CascadeMux I__779 (
            .O(N__9928),
            .I(N__9925));
    InMux I__778 (
            .O(N__9925),
            .I(N__9922));
    LocalMux I__777 (
            .O(N__9922),
            .I(\sb_translator_1.cnt_RNIKMBOZ0Z_9 ));
    CascadeMux I__776 (
            .O(N__9919),
            .I(N__9916));
    InMux I__775 (
            .O(N__9916),
            .I(N__9913));
    LocalMux I__774 (
            .O(N__9913),
            .I(\sb_translator_1.cnt_RNI6O3VZ0Z_10 ));
    InMux I__773 (
            .O(N__9910),
            .I(N__9907));
    LocalMux I__772 (
            .O(N__9907),
            .I(\sb_translator_1.cnt_RNIO5UPZ0Z_11 ));
    CascadeMux I__771 (
            .O(N__9904),
            .I(N__9901));
    InMux I__770 (
            .O(N__9901),
            .I(N__9898));
    LocalMux I__769 (
            .O(N__9898),
            .I(\sb_translator_1.cnt_RNISAVPZ0Z_12 ));
    CascadeMux I__768 (
            .O(N__9895),
            .I(N__9892));
    InMux I__767 (
            .O(N__9892),
            .I(N__9889));
    LocalMux I__766 (
            .O(N__9889),
            .I(\sb_translator_1.cnt_i_0 ));
    CascadeMux I__765 (
            .O(N__9886),
            .I(N__9883));
    InMux I__764 (
            .O(N__9883),
            .I(N__9880));
    LocalMux I__763 (
            .O(N__9880),
            .I(\sb_translator_1.cnt_i_1 ));
    CascadeMux I__762 (
            .O(N__9877),
            .I(N__9874));
    InMux I__761 (
            .O(N__9874),
            .I(N__9871));
    LocalMux I__760 (
            .O(N__9871),
            .I(\sb_translator_1.cnt_RNIOI3OZ0Z_2 ));
    InMux I__759 (
            .O(N__9868),
            .I(N__9865));
    LocalMux I__758 (
            .O(N__9865),
            .I(\sb_translator_1.cnt_RNISN4OZ0Z_3 ));
    INV \INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_1__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27512));
    INV \INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_2__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27519));
    INV \INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_10__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27462));
    INV \INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_5__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27430));
    INV \INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_11__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27477));
    INV \INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_0__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27446));
    INV \INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_4__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27423));
    INV \INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_6__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27442));
    INV \INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_3__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27419));
    INV \INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_13__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27504));
    INV \INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_12__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27491));
    INV \INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_7__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27456));
    INV \INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_8__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27472));
    INV \INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN  (
            .O(\INVgenblk1_genblk1_9__ram_i.mem_mem_0_0RCLKN_net ),
            .I(N__27487));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(\sb_translator_1.state56_a_5_cry_6 ),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(\sb_translator_1.state56_a_5_cry_14 ),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\ws2812.un6_data_cry_7 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\ws2812.un1_bit_counter_12_cry_7 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(\sb_translator_1.un1_num_leds_0_cry_8 ),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(\sb_translator_1.cnt_leds_cry_7 ),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\sb_translator_1.cnt_leds_cry_15 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(\sb_translator_1.cnt19_cry_7 ),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(\sb_translator_1.cnt19_cry_15 ),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(\sb_translator_1.cnt19_cry_25 ),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\sb_translator_1.cnt19_cry_33 ),
            .carryinitout(bfn_1_7_0_));
    ICE_GB \sb_translator_1.state_RNI6JH4_1  (
            .USERSIGNALTOGLOBALBUFFER(N__22798),
            .GLOBALBUFFEROUTPUT(\sb_translator_1.state_g_1 ));
    defparam OSCInst0.CLKHF_DIV="0b00";
    SB_HFOSC OSCInst0 (
            .CLKHFPU(N__26124),
            .CLKHFEN(N__26123),
            .CLKHF(clk_sb));
    ICE_GB \sb_translator_1.state_leds_RNIVONR_0  (
            .USERSIGNALTOGLOBALBUFFER(N__18010),
            .GLOBALBUFFEROUTPUT(\sb_translator_1.state_leds_2_sqmuxa_g ));
    ICE_GB reset_n_input_RNIVGR4_0 (
            .USERSIGNALTOGLOBALBUFFER(N__11245),
            .GLOBALBUFFEROUTPUT(reset_n_i_g));
    ICE_GB \spi_slave_1.bitcnt_rx_RNIPNM61_0_4  (
            .USERSIGNALTOGLOBALBUFFER(N__10069),
            .GLOBALBUFFEROUTPUT(\spi_slave_1.un3_mosi_data_out_g ));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \spi_slave_1.clk_RNIVAC01_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__10795),
            .GLOBALBUFFEROUTPUT(\spi_slave_1.bitcnt_rxe_0_i_g ));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \sb_translator_1.instr_tx_LC_0_10_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tx_LC_0_10_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tx_LC_0_10_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \sb_translator_1.instr_tx_LC_0_10_4  (
            .in0(N__23998),
            .in1(N__10761),
            .in2(_gnd_net_),
            .in3(N__22072),
            .lcout(miso_tx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27439),
            .ce(),
            .sr(N__27107));
    defparam \sb_translator_1.cnt_RNI4OM7_0_LC_1_3_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI4OM7_0_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI4OM7_0_LC_1_3_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \sb_translator_1.cnt_RNI4OM7_0_LC_1_3_0  (
            .in0(N__12513),
            .in1(N__19108),
            .in2(N__9895),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_i_0 ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\sb_translator_1.cnt19_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI1TPB_1_LC_1_3_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI1TPB_1_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI1TPB_1_LC_1_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI1TPB_1_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__11041),
            .in2(N__9886),
            .in3(N__12471),
            .lcout(\sb_translator_1.cnt_i_1 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_0 ),
            .carryout(\sb_translator_1.cnt19_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIOI3O_2_LC_1_3_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNIOI3O_2_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIOI3O_2_LC_1_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNIOI3O_2_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__11032),
            .in2(N__9877),
            .in3(N__12438),
            .lcout(\sb_translator_1.cnt_RNIOI3OZ0Z_2 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_1 ),
            .carryout(\sb_translator_1.cnt19_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNISN4O_3_LC_1_3_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNISN4O_3_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNISN4O_3_LC_1_3_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNISN4O_3_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__9868),
            .in2(N__11020),
            .in3(N__14628),
            .lcout(\sb_translator_1.cnt_RNISN4OZ0Z_3 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_2 ),
            .carryout(\sb_translator_1.cnt19_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI0T5O_4_LC_1_3_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI0T5O_4_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI0T5O_4_LC_1_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI0T5O_4_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__11005),
            .in2(N__9970),
            .in3(N__22560),
            .lcout(\sb_translator_1.cnt_RNI0T5OZ0Z_4 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_3 ),
            .carryout(\sb_translator_1.cnt19_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI427O_5_LC_1_3_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI427O_5_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI427O_5_LC_1_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI427O_5_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__10993),
            .in2(N__9961),
            .in3(N__14589),
            .lcout(\sb_translator_1.cnt_RNI427OZ0Z_5 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_4 ),
            .carryout(\sb_translator_1.cnt19_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI878O_6_LC_1_3_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI878O_6_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI878O_6_LC_1_3_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \sb_translator_1.cnt_RNI878O_6_LC_1_3_6  (
            .in0(N__22506),
            .in1(N__9952),
            .in2(N__10981),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_RNI878OZ0Z_6 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_5 ),
            .carryout(\sb_translator_1.cnt19_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNICC9O_7_LC_1_3_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNICC9O_7_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNICC9O_7_LC_1_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNICC9O_7_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(N__10966),
            .in2(N__9946),
            .in3(N__22927),
            .lcout(\sb_translator_1.cnt_RNICC9OZ0Z_7 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_6 ),
            .carryout(\sb_translator_1.cnt19_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIGHAO_8_LC_1_4_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNIGHAO_8_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIGHAO_8_LC_1_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNIGHAO_8_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__10954),
            .in2(N__9937),
            .in3(N__21446),
            .lcout(\sb_translator_1.cnt_RNIGHAOZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(\sb_translator_1.cnt19_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIKMBO_9_LC_1_4_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNIKMBO_9_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIKMBO_9_LC_1_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNIKMBO_9_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(N__11143),
            .in2(N__9928),
            .in3(N__10564),
            .lcout(\sb_translator_1.cnt_RNIKMBOZ0Z_9 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_8 ),
            .carryout(\sb_translator_1.cnt19_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI6O3V_10_LC_1_4_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI6O3V_10_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI6O3V_10_LC_1_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI6O3V_10_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(N__11131),
            .in2(N__9919),
            .in3(N__17291),
            .lcout(\sb_translator_1.cnt_RNI6O3VZ0Z_10 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_9 ),
            .carryout(\sb_translator_1.cnt19_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIO5UP_11_LC_1_4_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNIO5UP_11_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIO5UP_11_LC_1_4_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \sb_translator_1.cnt_RNIO5UP_11_LC_1_4_3  (
            .in0(N__17358),
            .in1(N__9910),
            .in2(N__11119),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_RNIO5UPZ0Z_11 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_10 ),
            .carryout(\sb_translator_1.cnt19_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNISAVP_12_LC_1_4_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNISAVP_12_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNISAVP_12_LC_1_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNISAVP_12_LC_1_4_4  (
            .in0(_gnd_net_),
            .in1(N__11104),
            .in2(N__9904),
            .in3(N__10531),
            .lcout(\sb_translator_1.cnt_RNISAVPZ0Z_12 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_11 ),
            .carryout(\sb_translator_1.cnt19_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI0G0Q_13_LC_1_4_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI0G0Q_13_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI0G0Q_13_LC_1_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI0G0Q_13_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(N__11092),
            .in2(N__10027),
            .in3(N__10423),
            .lcout(\sb_translator_1.cnt_RNI0G0QZ0Z_13 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_12 ),
            .carryout(\sb_translator_1.cnt19_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI4L1Q_14_LC_1_4_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI4L1Q_14_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI4L1Q_14_LC_1_4_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \sb_translator_1.cnt_RNI4L1Q_14_LC_1_4_6  (
            .in0(N__10402),
            .in1(N__11080),
            .in2(N__10015),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_RNI4L1QZ0Z_14 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_13 ),
            .carryout(\sb_translator_1.cnt19_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNI8Q2Q_15_LC_1_4_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNI8Q2Q_15_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNI8Q2Q_15_LC_1_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNI8Q2Q_15_LC_1_4_7  (
            .in0(_gnd_net_),
            .in1(N__11068),
            .in2(N__10003),
            .in3(N__10381),
            .lcout(\sb_translator_1.cnt_RNI8Q2QZ0Z_15 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_14 ),
            .carryout(\sb_translator_1.cnt19_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIQ4UI_16_LC_1_5_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNIQ4UI_16_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIQ4UI_16_LC_1_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_RNIQ4UI_16_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__11053),
            .in2(N__9991),
            .in3(N__10359),
            .lcout(\sb_translator_1.cnt_i_16 ),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\sb_translator_1.cnt19_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNIOCIR9_5_LC_1_5_1 .C_ON=1'b1;
    defparam \sb_translator_1.state_RNIOCIR9_5_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIOCIR9_5_LC_1_5_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \sb_translator_1.state_RNIOCIR9_5_LC_1_5_1  (
            .in0(N__10281),
            .in1(N__23011),
            .in2(_gnd_net_),
            .in3(N__9982),
            .lcout(\sb_translator_1.state_RNIOCIR9Z0Z_5 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_16 ),
            .carryout(\sb_translator_1.cnt19_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt19_cry_18_THRU_LUT4_0_LC_1_5_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt19_cry_18_THRU_LUT4_0_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt19_cry_18_THRU_LUT4_0_LC_1_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.cnt19_cry_18_THRU_LUT4_0_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__12508),
            .in2(_gnd_net_),
            .in3(N__9979),
            .lcout(\sb_translator_1.cnt19_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_18 ),
            .carryout(\sb_translator_1.cnt19_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_1_LC_1_5_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_1_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_1_LC_1_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_1_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__12461),
            .in2(_gnd_net_),
            .in3(N__9976),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_20 ),
            .carryout(\sb_translator_1.cnt19_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_2_LC_1_5_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_2_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_2_LC_1_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_2_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__12434),
            .in2(_gnd_net_),
            .in3(N__9973),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_21 ),
            .carryout(\sb_translator_1.cnt19_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_3_LC_1_5_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_3_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_3_LC_1_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_3_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__14624),
            .in2(_gnd_net_),
            .in3(N__10054),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_22 ),
            .carryout(\sb_translator_1.cnt19_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_4_LC_1_5_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_4_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_4_LC_1_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_4_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(N__22556),
            .in2(_gnd_net_),
            .in3(N__10051),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_23 ),
            .carryout(\sb_translator_1.cnt19_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_5_LC_1_5_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_5_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_5_LC_1_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_5_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__14585),
            .in2(_gnd_net_),
            .in3(N__10048),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_24 ),
            .carryout(\sb_translator_1.cnt19_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_6_LC_1_6_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_6_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_6_LC_1_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_6_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__22502),
            .in2(_gnd_net_),
            .in3(N__10045),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\sb_translator_1.cnt19_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_7_LC_1_6_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_7_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_7_LC_1_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_7_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__22919),
            .in2(_gnd_net_),
            .in3(N__10042),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_26 ),
            .carryout(\sb_translator_1.cnt19_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_8_LC_1_6_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_8_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_8_LC_1_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_8_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__21447),
            .in2(_gnd_net_),
            .in3(N__10039),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_27 ),
            .carryout(\sb_translator_1.cnt19_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_9_LC_1_6_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_9_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_9_LC_1_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_9_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__10556),
            .in2(_gnd_net_),
            .in3(N__10036),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_28 ),
            .carryout(\sb_translator_1.cnt19_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_10_LC_1_6_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_10_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_10_LC_1_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_10_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__17292),
            .in2(_gnd_net_),
            .in3(N__10033),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_29 ),
            .carryout(\sb_translator_1.cnt19_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_11_LC_1_6_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_11_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_11_LC_1_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_11_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__17346),
            .in2(_gnd_net_),
            .in3(N__10030),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_30 ),
            .carryout(\sb_translator_1.cnt19_cry_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_12_LC_1_6_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_12_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_12_LC_1_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_12_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__10517),
            .in2(_gnd_net_),
            .in3(N__10084),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_31 ),
            .carryout(\sb_translator_1.cnt19_cry_32 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_13_LC_1_6_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_13_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_13_LC_1_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_13_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__10422),
            .in2(_gnd_net_),
            .in3(N__10081),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_32 ),
            .carryout(\sb_translator_1.cnt19_cry_33 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_14_LC_1_7_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_14_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_14_LC_1_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_14_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__10401),
            .in2(_gnd_net_),
            .in3(N__10078),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\sb_translator_1.cnt19_cry_34 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_15_LC_1_7_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_RNO_0_15_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_15_LC_1_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_15_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__10380),
            .in2(_gnd_net_),
            .in3(N__10075),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt19_cry_34 ),
            .carryout(\sb_translator_1.cnt19_cry_35 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNO_0_16_LC_1_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNO_0_16_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_16_LC_1_7_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \sb_translator_1.cnt_RNO_0_16_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__10360),
            .in2(_gnd_net_),
            .in3(N__10072),
            .lcout(\sb_translator_1.cnt_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNIKJOC_5_LC_1_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIKJOC_5_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIKJOC_5_LC_1_7_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \sb_translator_1.state_RNIKJOC_5_LC_1_7_4  (
            .in0(N__10282),
            .in1(N__22066),
            .in2(_gnd_net_),
            .in3(N__16853),
            .lcout(\sb_translator_1.state_RNIKJOCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_tmp_23_LC_1_8_2 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_23_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_23_LC_1_8_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_23_LC_1_8_2  (
            .in0(N__16844),
            .in1(N__22762),
            .in2(N__10615),
            .in3(N__22071),
            .lcout(\sb_translator_1.instr_tmpZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27434),
            .ce(),
            .sr(N__27088));
    defparam \sb_translator_1.instr_tmp_21_LC_1_8_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_21_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_21_LC_1_8_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \sb_translator_1.instr_tmp_21_LC_1_8_4  (
            .in0(N__16843),
            .in1(N__22070),
            .in2(N__10447),
            .in3(N__22644),
            .lcout(\sb_translator_1.instr_tmpZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27434),
            .ce(),
            .sr(N__27088));
    defparam \sb_translator_1.instr_tmp_18_LC_1_8_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_18_LC_1_8_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_18_LC_1_8_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_18_LC_1_8_5  (
            .in0(N__17680),
            .in1(N__22073),
            .in2(N__10492),
            .in3(N__16842),
            .lcout(\sb_translator_1.instr_tmpZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27434),
            .ce(),
            .sr(N__27088));
    defparam \spi_slave_1.bitcnt_rx_RNIPNM61_4_LC_1_9_0 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_rx_RNIPNM61_4_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_rx_RNIPNM61_4_LC_1_9_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \spi_slave_1.bitcnt_rx_RNIPNM61_4_LC_1_9_0  (
            .in0(N__10172),
            .in1(N__10141),
            .in2(_gnd_net_),
            .in3(N__10130),
            .lcout(\spi_slave_1.bitcnt_rx_RNIPNM61Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_rx_RNI3EGR_1_LC_1_9_1 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_rx_RNI3EGR_1_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_rx_RNI3EGR_1_LC_1_9_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \spi_slave_1.bitcnt_rx_RNI3EGR_1_LC_1_9_1  (
            .in0(N__10191),
            .in1(N__10098),
            .in2(N__11876),
            .in3(N__10113),
            .lcout(\spi_slave_1.un3_mosi_data_out_3 ),
            .ltout(\spi_slave_1.un3_mosi_data_out_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.mosi_rx_LC_1_9_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_rx_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_rx_LC_1_9_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \spi_slave_1.mosi_rx_LC_1_9_2  (
            .in0(N__10173),
            .in1(_gnd_net_),
            .in2(N__10135),
            .in3(N__10131),
            .lcout(mosi_rx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27440),
            .ce(),
            .sr(N__27095));
    defparam \sb_translator_1.instr_tmp_19_LC_1_9_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_19_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_19_LC_1_9_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_19_LC_1_9_4  (
            .in0(N__22064),
            .in1(N__17623),
            .in2(N__10477),
            .in3(N__16826),
            .lcout(\sb_translator_1.instr_tmpZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27440),
            .ce(),
            .sr(N__27095));
    defparam \sb_translator_1.instr_tmp_20_LC_1_9_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_20_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_20_LC_1_9_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_20_LC_1_9_5  (
            .in0(N__16827),
            .in1(N__17572),
            .in2(N__10462),
            .in3(N__22065),
            .lcout(\sb_translator_1.instr_tmpZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27440),
            .ce(),
            .sr(N__27095));
    defparam \sb_translator_1.state_RNIH20C_0_LC_1_9_6 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIH20C_0_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIH20C_0_LC_1_9_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \sb_translator_1.state_RNIH20C_0_LC_1_9_6  (
            .in0(N__22063),
            .in1(N__16825),
            .in2(_gnd_net_),
            .in3(N__22643),
            .lcout(\sb_translator_1.N_1087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_6_0_0_a2_1_9_LC_1_9_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_1_9_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_1_9_LC_1_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \sb_translator_1.ram_sel_6_0_0_a2_1_9_LC_1_9_7  (
            .in0(N__17622),
            .in1(N__17571),
            .in2(_gnd_net_),
            .in3(N__17679),
            .lcout(\sb_translator_1.ram_sel_6_0_0_a2_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_rx_0_LC_1_10_0 .C_ON=1'b1;
    defparam \spi_slave_1.bitcnt_rx_0_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.bitcnt_rx_0_LC_1_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_rx_0_LC_1_10_0  (
            .in0(N__10702),
            .in1(N__10132),
            .in2(_gnd_net_),
            .in3(N__10117),
            .lcout(\spi_slave_1.bitcnt_rxZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\spi_slave_1.bitcnt_rx_cry_0 ),
            .clk(N__27448),
            .ce(N__12064),
            .sr(N__27100));
    defparam \spi_slave_1.bitcnt_rx_1_LC_1_10_1 .C_ON=1'b1;
    defparam \spi_slave_1.bitcnt_rx_1_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.bitcnt_rx_1_LC_1_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_rx_1_LC_1_10_1  (
            .in0(N__10710),
            .in1(N__10114),
            .in2(_gnd_net_),
            .in3(N__10102),
            .lcout(\spi_slave_1.bitcnt_rxZ0Z_1 ),
            .ltout(),
            .carryin(\spi_slave_1.bitcnt_rx_cry_0 ),
            .carryout(\spi_slave_1.bitcnt_rx_cry_1 ),
            .clk(N__27448),
            .ce(N__12064),
            .sr(N__27100));
    defparam \spi_slave_1.bitcnt_rx_2_LC_1_10_2 .C_ON=1'b1;
    defparam \spi_slave_1.bitcnt_rx_2_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.bitcnt_rx_2_LC_1_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_rx_2_LC_1_10_2  (
            .in0(N__10703),
            .in1(N__10099),
            .in2(_gnd_net_),
            .in3(N__10087),
            .lcout(\spi_slave_1.bitcnt_rxZ0Z_2 ),
            .ltout(),
            .carryin(\spi_slave_1.bitcnt_rx_cry_1 ),
            .carryout(\spi_slave_1.bitcnt_rx_cry_2 ),
            .clk(N__27448),
            .ce(N__12064),
            .sr(N__27100));
    defparam \spi_slave_1.bitcnt_rx_3_LC_1_10_3 .C_ON=1'b1;
    defparam \spi_slave_1.bitcnt_rx_3_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.bitcnt_rx_3_LC_1_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_rx_3_LC_1_10_3  (
            .in0(N__10711),
            .in1(N__10192),
            .in2(_gnd_net_),
            .in3(N__10180),
            .lcout(\spi_slave_1.bitcnt_rxZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_1.bitcnt_rx_cry_2 ),
            .carryout(\spi_slave_1.bitcnt_rx_cry_3 ),
            .clk(N__27448),
            .ce(N__12064),
            .sr(N__27100));
    defparam \spi_slave_1.bitcnt_rx_4_LC_1_10_4 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_rx_4_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.bitcnt_rx_4_LC_1_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_rx_4_LC_1_10_4  (
            .in0(N__10704),
            .in1(N__10174),
            .in2(_gnd_net_),
            .in3(N__10177),
            .lcout(\spi_slave_1.bitcnt_rxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27448),
            .ce(N__12064),
            .sr(N__27100));
    defparam \spi_slave_1.miso_en_LC_1_11_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_en_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_en_LC_1_11_1 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \spi_slave_1.miso_en_LC_1_11_1  (
            .in0(N__10159),
            .in1(N__10885),
            .in2(N__11877),
            .in3(N__10861),
            .lcout(miso_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27454),
            .ce(),
            .sr(N__27110));
    defparam \sb_translator_1.instr_tmp_17_LC_1_11_6 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_17_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_17_LC_1_11_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_17_LC_1_11_6  (
            .in0(N__11335),
            .in1(N__22075),
            .in2(N__14667),
            .in3(N__16852),
            .lcout(\sb_translator_1.instr_tmpZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27454),
            .ce(),
            .sr(N__27110));
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_c_LC_1_12_0 .C_ON=1'b1;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_slave_1.un1_bitcnt_tx_1_cry_0_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__18512),
            .in2(N__10783),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\spi_slave_1.un1_bitcnt_tx_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_LUT4_0_LC_1_12_1 .C_ON=1'b1;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_LUT4_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_LUT4_0_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_LUT4_0_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__11941),
            .in2(_gnd_net_),
            .in3(N__10153),
            .lcout(\spi_slave_1.un1_bitcnt_tx_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_1.un1_bitcnt_tx_1_cry_0 ),
            .carryout(\spi_slave_1.un1_bitcnt_tx_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_LUT4_0_LC_1_12_2 .C_ON=1'b1;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_LUT4_0_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_LUT4_0_LC_1_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_LUT4_0_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__11694),
            .in2(_gnd_net_),
            .in3(N__10150),
            .lcout(\spi_slave_1.un1_bitcnt_tx_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_1.un1_bitcnt_tx_1_cry_1 ),
            .carryout(\spi_slave_1.un1_bitcnt_tx_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_3_LC_1_12_3 .C_ON=1'b1;
    defparam \spi_slave_1.bitcnt_tx_3_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.bitcnt_tx_3_LC_1_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_1.bitcnt_tx_3_LC_1_12_3  (
            .in0(N__27159),
            .in1(N__10860),
            .in2(_gnd_net_),
            .in3(N__10147),
            .lcout(\spi_slave_1.bitcnt_txZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_1.un1_bitcnt_tx_1_cry_2 ),
            .carryout(\spi_slave_1.un1_bitcnt_tx_1_cry_3 ),
            .clk(N__27464),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_4_LC_1_12_4 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_4_LC_1_12_4 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.bitcnt_tx_4_LC_1_12_4 .LUT_INIT=16'b1010101110111010;
    LogicCell40 \spi_slave_1.bitcnt_tx_4_LC_1_12_4  (
            .in0(N__27158),
            .in1(N__10914),
            .in2(N__18580),
            .in3(N__10144),
            .lcout(\spi_slave_1.bitcnt_txZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27464),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_2_LC_1_12_5 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_2_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.bitcnt_tx_2_LC_1_12_5 .LUT_INIT=16'b1100110111001110;
    LogicCell40 \spi_slave_1.bitcnt_tx_2_LC_1_12_5  (
            .in0(N__11695),
            .in1(N__27157),
            .in2(N__10921),
            .in3(N__10204),
            .lcout(\spi_slave_1.bitcnt_txZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27464),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_1_LC_1_12_6 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_1_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.bitcnt_tx_1_LC_1_12_6 .LUT_INIT=16'b1111000111110010;
    LogicCell40 \spi_slave_1.bitcnt_tx_1_LC_1_12_6  (
            .in0(N__11942),
            .in1(N__10915),
            .in2(N__27160),
            .in3(N__10198),
            .lcout(\spi_slave_1.bitcnt_txZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27464),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_2_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_2_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_2_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_2_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.mosi_data_in_18_LC_2_3_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_18_LC_2_3_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_18_LC_2_3_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_18_LC_2_3_0  (
            .in0(N__12087),
            .in1(N__12186),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_19_LC_2_3_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_19_LC_2_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_19_LC_2_3_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_19_LC_2_3_1  (
            .in0(N__12324),
            .in1(_gnd_net_),
            .in2(N__12224),
            .in3(N__10263),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_20_LC_2_3_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_20_LC_2_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_20_LC_2_3_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_20_LC_2_3_2  (
            .in0(N__10251),
            .in1(N__12190),
            .in2(_gnd_net_),
            .in3(N__12325),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_21_LC_2_3_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_21_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_21_LC_2_3_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_21_LC_2_3_3  (
            .in0(N__12326),
            .in1(_gnd_net_),
            .in2(N__12225),
            .in3(N__10239),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_22_LC_2_3_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_22_LC_2_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_22_LC_2_3_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_22_LC_2_3_4  (
            .in0(N__10227),
            .in1(N__12194),
            .in2(_gnd_net_),
            .in3(N__12327),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_23_LC_2_3_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_23_LC_2_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_23_LC_2_3_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_23_LC_2_3_5  (
            .in0(N__12328),
            .in1(_gnd_net_),
            .in2(N__12226),
            .in3(N__10215),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_8_LC_2_3_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_8_LC_2_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_8_LC_2_3_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_8_LC_2_3_6  (
            .in0(N__13198),
            .in1(N__12198),
            .in2(_gnd_net_),
            .in3(N__12329),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_in_9_LC_2_3_7 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_9_LC_2_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_9_LC_2_3_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_9_LC_2_3_7  (
            .in0(N__12330),
            .in1(_gnd_net_),
            .in2(N__12227),
            .in3(N__12015),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27421),
            .ce(N__12062),
            .sr(N__27065));
    defparam \spi_slave_1.mosi_data_out_17_LC_2_4_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_17_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_17_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_17_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12088),
            .lcout(mosi_data_out_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_23_LC_2_4_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_23_LC_2_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_23_LC_2_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_23_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10270),
            .lcout(mosi_data_out_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_18_LC_2_4_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_18_LC_2_4_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_18_LC_2_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_18_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10264),
            .lcout(mosi_data_out_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_19_LC_2_4_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_19_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_19_LC_2_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_19_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10252),
            .lcout(mosi_data_out_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_1_LC_2_4_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_1_LC_2_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_1_LC_2_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_1.mosi_data_out_1_LC_2_4_4  (
            .in0(N__11161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(mosi_data_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_20_LC_2_4_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_20_LC_2_4_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_20_LC_2_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_20_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10240),
            .lcout(mosi_data_out_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_21_LC_2_4_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_21_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_21_LC_2_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_21_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10228),
            .lcout(mosi_data_out_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \spi_slave_1.mosi_data_out_22_LC_2_4_7 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_22_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_22_LC_2_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_22_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10216),
            .lcout(mosi_data_out_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27422),
            .ce(N__18424),
            .sr(N__27067));
    defparam \sb_translator_1.cnt_10_LC_2_5_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_10_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_10_LC_2_5_0 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_10_LC_2_5_0  (
            .in0(N__22763),
            .in1(N__17094),
            .in2(N__17220),
            .in3(N__10330),
            .lcout(\sb_translator_1.cntZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_2_LC_2_5_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_2_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_2_LC_2_5_1 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_2_LC_2_5_1  (
            .in0(N__17090),
            .in1(N__17177),
            .in2(N__22786),
            .in3(N__10324),
            .lcout(\sb_translator_1.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_3_LC_2_5_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_3_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_3_LC_2_5_2 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_3_LC_2_5_2  (
            .in0(N__22764),
            .in1(N__17095),
            .in2(N__17221),
            .in3(N__10318),
            .lcout(\sb_translator_1.cntZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_4_LC_2_5_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_4_LC_2_5_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_4_LC_2_5_3 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_4_LC_2_5_3  (
            .in0(N__17091),
            .in1(N__17178),
            .in2(N__22787),
            .in3(N__10312),
            .lcout(\sb_translator_1.cntZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_5_LC_2_5_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_5_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_5_LC_2_5_4 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_5_LC_2_5_4  (
            .in0(N__22765),
            .in1(N__17096),
            .in2(N__17222),
            .in3(N__10306),
            .lcout(\sb_translator_1.cntZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_6_LC_2_5_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_6_LC_2_5_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_6_LC_2_5_5 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_6_LC_2_5_5  (
            .in0(N__17092),
            .in1(N__17179),
            .in2(N__22788),
            .in3(N__10300),
            .lcout(\sb_translator_1.cntZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_7_LC_2_5_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_7_LC_2_5_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_7_LC_2_5_6 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_7_LC_2_5_6  (
            .in0(N__22766),
            .in1(N__17097),
            .in2(N__17223),
            .in3(N__10294),
            .lcout(\sb_translator_1.cntZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.cnt_8_LC_2_5_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_8_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_8_LC_2_5_7 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_8_LC_2_5_7  (
            .in0(N__17093),
            .in1(N__17180),
            .in2(N__22789),
            .in3(N__10288),
            .lcout(\sb_translator_1.cntZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27427),
            .ce(),
            .sr(N__27070));
    defparam \sb_translator_1.state_5_LC_2_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.state_5_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.state_5_LC_2_6_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \sb_translator_1.state_5_LC_2_6_0  (
            .in0(N__17199),
            .in1(N__22735),
            .in2(_gnd_net_),
            .in3(N__17104),
            .lcout(\sb_translator_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_RNO_0_0_LC_2_6_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNO_0_0_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNO_0_0_LC_2_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \sb_translator_1.cnt_RNO_0_0_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__12512),
            .in2(_gnd_net_),
            .in3(N__16881),
            .lcout(),
            .ltout(\sb_translator_1.cnt_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_0_LC_2_6_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_0_LC_2_6_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_0_LC_2_6_2 .LUT_INIT=16'b1001000011110000;
    LogicCell40 \sb_translator_1.cnt_0_LC_2_6_2  (
            .in0(N__17196),
            .in1(N__22734),
            .in2(N__10432),
            .in3(N__17103),
            .lcout(\sb_translator_1.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_13_LC_2_6_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_13_LC_2_6_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_13_LC_2_6_3 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_13_LC_2_6_3  (
            .in0(N__17098),
            .in1(N__17200),
            .in2(N__22779),
            .in3(N__10429),
            .lcout(\sb_translator_1.cntZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_14_LC_2_6_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_14_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_14_LC_2_6_4 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_14_LC_2_6_4  (
            .in0(N__17197),
            .in1(N__17101),
            .in2(N__22782),
            .in3(N__10408),
            .lcout(\sb_translator_1.cntZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_15_LC_2_6_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_15_LC_2_6_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_15_LC_2_6_5 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_15_LC_2_6_5  (
            .in0(N__17099),
            .in1(N__17201),
            .in2(N__22780),
            .in3(N__10387),
            .lcout(\sb_translator_1.cntZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_16_LC_2_6_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_16_LC_2_6_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_16_LC_2_6_6 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_16_LC_2_6_6  (
            .in0(N__17198),
            .in1(N__17102),
            .in2(N__22783),
            .in3(N__10366),
            .lcout(\sb_translator_1.cntZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_1_LC_2_6_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_1_LC_2_6_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_1_LC_2_6_7 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_1_LC_2_6_7  (
            .in0(N__17100),
            .in1(N__17202),
            .in2(N__22781),
            .in3(N__10348),
            .lcout(\sb_translator_1.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27429),
            .ce(),
            .sr(N__27074));
    defparam \sb_translator_1.cnt_11_LC_2_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_11_LC_2_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_11_LC_2_7_0 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_11_LC_2_7_0  (
            .in0(N__17105),
            .in1(N__22760),
            .in2(N__17227),
            .in3(N__10342),
            .lcout(\sb_translator_1.cntZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27435),
            .ce(),
            .sr(N__27077));
    defparam \sb_translator_1.cnt_12_LC_2_7_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_12_LC_2_7_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_12_LC_2_7_1 .LUT_INIT=16'b1011011100000000;
    LogicCell40 \sb_translator_1.cnt_12_LC_2_7_1  (
            .in0(N__22759),
            .in1(N__17107),
            .in2(N__17234),
            .in3(N__10336),
            .lcout(\sb_translator_1.cntZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27435),
            .ce(),
            .sr(N__27077));
    defparam \sb_translator_1.cnt_9_LC_2_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_9_LC_2_7_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_9_LC_2_7_2 .LUT_INIT=16'b1101011100000000;
    LogicCell40 \sb_translator_1.cnt_9_LC_2_7_2  (
            .in0(N__17106),
            .in1(N__22761),
            .in2(N__17228),
            .in3(N__10570),
            .lcout(\sb_translator_1.cntZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27435),
            .ce(),
            .sr(N__27077));
    defparam \sb_translator_1.cnt_RNIJ7EF_1_9_LC_2_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNIJ7EF_1_9_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIJ7EF_1_9_LC_2_7_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \sb_translator_1.cnt_RNIJ7EF_1_9_LC_2_7_3  (
            .in0(N__22057),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__10557),
            .lcout(\sb_translator_1.cnt_RNIJ7EF_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIJ7EF_2_9_LC_2_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNIJ7EF_2_9_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIJ7EF_2_9_LC_2_7_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \sb_translator_1.cnt_RNIJ7EF_2_9_LC_2_7_4  (
            .in0(N__10558),
            .in1(_gnd_net_),
            .in2(N__10529),
            .in3(N__22059),
            .lcout(\sb_translator_1.cnt_RNIJ7EF_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIJ7EF_0_9_LC_2_7_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNIJ7EF_0_9_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIJ7EF_0_9_LC_2_7_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \sb_translator_1.cnt_RNIJ7EF_0_9_LC_2_7_5  (
            .in0(N__22058),
            .in1(N__10522),
            .in2(_gnd_net_),
            .in3(N__10559),
            .lcout(\sb_translator_1.N_1088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNIJ7EF_9_LC_2_7_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNIJ7EF_9_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNIJ7EF_9_LC_2_7_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \sb_translator_1.cnt_RNIJ7EF_9_LC_2_7_6  (
            .in0(N__10560),
            .in1(_gnd_net_),
            .in2(N__10530),
            .in3(N__22060),
            .lcout(\sb_translator_1.N_1092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_tmp_22_LC_2_7_7 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_22_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_22_LC_2_7_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \sb_translator_1.instr_tmp_22_LC_2_7_7  (
            .in0(N__22061),
            .in1(N__17203),
            .in2(N__10630),
            .in3(N__16864),
            .lcout(\sb_translator_1.instr_tmpZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27435),
            .ce(),
            .sr(N__27077));
    defparam \sb_translator_1.instr_out_18_LC_2_8_0 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_18_LC_2_8_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_18_LC_2_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_18_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10491),
            .lcout(miso_data_in_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_19_LC_2_8_1 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_19_LC_2_8_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_19_LC_2_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_19_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10476),
            .lcout(miso_data_in_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_20_LC_2_8_2 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_20_LC_2_8_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_20_LC_2_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.instr_out_20_LC_2_8_2  (
            .in0(N__10461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(miso_data_in_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_21_LC_2_8_3 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_21_LC_2_8_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_21_LC_2_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_21_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10446),
            .lcout(miso_data_in_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_22_LC_2_8_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_22_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_22_LC_2_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_22_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10629),
            .lcout(miso_data_in_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_23_LC_2_8_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_23_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_23_LC_2_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_23_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10614),
            .lcout(miso_data_in_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_8_LC_2_8_6 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_8_LC_2_8_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_8_LC_2_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_8_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15621),
            .lcout(miso_data_in_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \sb_translator_1.instr_out_9_LC_2_8_7 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_9_LC_2_8_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_9_LC_2_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.instr_out_9_LC_2_8_7  (
            .in0(N__15408),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(miso_data_in_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27441),
            .ce(N__23993),
            .sr(N__27082));
    defparam \spi_slave_1.miso_data_out_19_LC_2_9_0 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_19_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_19_LC_2_9_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_slave_1.miso_data_out_19_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.miso_data_outZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_20_LC_2_9_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_20_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_20_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_20_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10594),
            .lcout(\spi_slave_1.miso_data_outZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_21_LC_2_9_2 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_21_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_21_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_21_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10588),
            .lcout(\spi_slave_1.miso_data_outZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_22_LC_2_9_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_22_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_22_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_22_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10582),
            .lcout(\spi_slave_1.miso_data_outZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_23_LC_2_9_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_23_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_23_LC_2_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_23_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10576),
            .lcout(\spi_slave_1.miso_data_outZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_5_LC_2_9_5 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_5_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_5_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_5_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24277),
            .lcout(\spi_slave_1.miso_data_outZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_8_LC_2_9_6 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_8_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_8_LC_2_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_8_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10717),
            .lcout(\spi_slave_1.miso_data_outZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_4_LC_2_9_7 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_4_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_4_LC_2_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_4_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24013),
            .lcout(\spi_slave_1.miso_data_outZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27449),
            .ce(N__14547),
            .sr(_gnd_net_));
    defparam \spi_slave_1.clk_RNIDBLL_1_LC_2_10_0 .C_ON=1'b0;
    defparam \spi_slave_1.clk_RNIDBLL_1_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.clk_RNIDBLL_1_LC_2_10_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \spi_slave_1.clk_RNIDBLL_1_LC_2_10_0  (
            .in0(N__12277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12146),
            .lcout(\spi_slave_1.clk_pos_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_18_LC_2_10_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_18_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_18_LC_2_10_1 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \spi_slave_1.miso_RNO_18_LC_2_10_1  (
            .in0(N__11524),
            .in1(N__18582),
            .in2(N__10687),
            .in3(N__18504),
            .lcout(),
            .ltout(\spi_slave_1.m81_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_16_LC_2_10_2 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_16_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_16_LC_2_10_2 .LUT_INIT=16'b0111000001111010;
    LogicCell40 \spi_slave_1.miso_RNO_16_LC_2_10_2  (
            .in0(N__18506),
            .in1(N__10678),
            .in2(N__10672),
            .in3(N__10669),
            .lcout(\spi_slave_1.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_15_LC_2_10_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_15_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_15_LC_2_10_3 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \spi_slave_1.miso_RNO_15_LC_2_10_3  (
            .in0(N__10663),
            .in1(N__18583),
            .in2(N__10657),
            .in3(N__18505),
            .lcout(),
            .ltout(\spi_slave_1.m60_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_10_LC_2_10_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_10_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_10_LC_2_10_4 .LUT_INIT=16'b0111000001111010;
    LogicCell40 \spi_slave_1.miso_RNO_10_LC_2_10_4  (
            .in0(N__18507),
            .in1(N__10648),
            .in2(N__10642),
            .in3(N__11770),
            .lcout(\spi_slave_1.miso_RNOZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.clk_0_LC_2_11_0 .C_ON=1'b0;
    defparam \spi_slave_1.clk_0_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.clk_0_LC_2_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_1.clk_0_LC_2_11_0  (
            .in0(N__10639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.clkZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27465),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.clk_RNIFQ8K3_1_LC_2_11_1 .C_ON=1'b0;
    defparam \spi_slave_1.clk_RNIFQ8K3_1_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.clk_RNIFQ8K3_1_LC_2_11_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \spi_slave_1.clk_RNIFQ8K3_1_LC_2_11_1  (
            .in0(N__12111),
            .in1(N__12267),
            .in2(N__11864),
            .in3(N__10830),
            .lcout(\spi_slave_1.bitcnt_tx10 ),
            .ltout(\spi_slave_1.bitcnt_tx10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_0_LC_2_11_2 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_0_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.bitcnt_tx_0_LC_2_11_2 .LUT_INIT=16'b1100110011011110;
    LogicCell40 \spi_slave_1.bitcnt_tx_0_LC_2_11_2  (
            .in0(N__18510),
            .in1(N__27153),
            .in2(N__10774),
            .in3(N__10919),
            .lcout(\spi_slave_1.bitcnt_txZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27465),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_2_LC_2_11_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_2_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_2_LC_2_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.miso_RNO_2_LC_2_11_3  (
            .in0(N__12112),
            .in1(N__12268),
            .in2(_gnd_net_),
            .in3(N__10831),
            .lcout(\spi_slave_1.N_96_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_7_LC_2_11_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_7_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_7_LC_2_11_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \spi_slave_1.miso_RNO_7_LC_2_11_4  (
            .in0(N__18509),
            .in1(N__10771),
            .in2(_gnd_net_),
            .in3(N__11758),
            .lcout(\spi_slave_1.miso_RNOZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.clk_1_LC_2_11_5 .C_ON=1'b0;
    defparam \spi_slave_1.clk_1_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.clk_1_LC_2_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_slave_1.clk_1_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__12269),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.clkZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27465),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_RNIQORT2_3_LC_2_11_6 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_RNIQORT2_3_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_tx_RNIQORT2_3_LC_2_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \spi_slave_1.bitcnt_tx_RNIQORT2_3_LC_2_11_6  (
            .in0(N__10883),
            .in1(N__10762),
            .in2(N__11863),
            .in3(N__10859),
            .lcout(\spi_slave_1.miso_data_out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_17_LC_2_11_7 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_17_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_17_LC_2_11_7 .LUT_INIT=16'b0011111101000100;
    LogicCell40 \spi_slave_1.miso_RNO_17_LC_2_11_7  (
            .in0(N__11512),
            .in1(N__18508),
            .in2(N__14566),
            .in3(N__11722),
            .lcout(\spi_slave_1.miso_RNOZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_11_LC_2_12_0 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_11_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_11_LC_2_12_0 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \spi_slave_1.miso_RNO_11_LC_2_12_0  (
            .in0(N__11934),
            .in1(N__10744),
            .in2(N__11697),
            .in3(N__10735),
            .lcout(),
            .ltout(\spi_slave_1.m48_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_5_LC_2_12_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_5_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_5_LC_2_12_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \spi_slave_1.miso_RNO_5_LC_2_12_1  (
            .in0(N__18454),
            .in1(N__10729),
            .in2(N__10720),
            .in3(N__11935),
            .lcout(),
            .ltout(\spi_slave_1.N_49_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_3_LC_2_12_2 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_3_LC_2_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \spi_slave_1.miso_RNO_3_LC_2_12_2  (
            .in0(N__10863),
            .in1(_gnd_net_),
            .in2(N__10939),
            .in3(N__11896),
            .lcout(),
            .ltout(\spi_slave_1.N_25_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_1_LC_2_12_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_1_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_1_LC_2_12_3 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \spi_slave_1.miso_RNO_1_LC_2_12_3  (
            .in0(N__11841),
            .in1(_gnd_net_),
            .in2(N__10936),
            .in3(N__10933),
            .lcout(\spi_slave_1.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_RNIP9N23_3_LC_2_12_4 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_RNIP9N23_3_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_tx_RNIP9N23_3_LC_2_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \spi_slave_1.bitcnt_tx_RNIP9N23_3_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__11274),
            .in2(_gnd_net_),
            .in3(N__10920),
            .lcout(\spi_slave_1.bitcnt_tx_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_0_LC_2_12_5 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_0_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_0_LC_2_12_5 .LUT_INIT=16'b0010000000101111;
    LogicCell40 \spi_slave_1.miso_RNO_0_LC_2_12_5  (
            .in0(N__10884),
            .in1(N__10864),
            .in2(N__11862),
            .in3(N__10891),
            .lcout(\spi_slave_1.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_RNIJITN1_2_LC_2_12_6 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_RNIJITN1_2_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_tx_RNIJITN1_2_LC_2_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \spi_slave_1.bitcnt_tx_RNIJITN1_2_LC_2_12_6  (
            .in0(N__11933),
            .in1(N__18563),
            .in2(N__11696),
            .in3(N__18511),
            .lcout(\spi_slave_1.N_94_mux ),
            .ltout(\spi_slave_1.N_94_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.bitcnt_tx_RNIGFSJ2_3_LC_2_12_7 .C_ON=1'b0;
    defparam \spi_slave_1.bitcnt_tx_RNIGFSJ2_3_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.bitcnt_tx_RNIGFSJ2_3_LC_2_12_7 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \spi_slave_1.bitcnt_tx_RNIGFSJ2_3_LC_2_12_7  (
            .in0(N__18564),
            .in1(_gnd_net_),
            .in2(N__10867),
            .in3(N__10862),
            .lcout(\spi_slave_1.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_LC_2_13_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_LC_2_13_1 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_LC_2_13_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \spi_slave_1.miso_LC_2_13_1  (
            .in0(N__10806),
            .in1(N__10822),
            .in2(_gnd_net_),
            .in3(N__10816),
            .lcout(miso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27480),
            .ce(),
            .sr(N__27113));
    defparam \spi_slave_1.clk_RNIVAC01_1_LC_4_1_7 .C_ON=1'b0;
    defparam \spi_slave_1.clk_RNIVAC01_1_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.clk_RNIVAC01_1_LC_4_1_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \spi_slave_1.clk_RNIVAC01_1_LC_4_1_7  (
            .in0(N__12202),
            .in1(N__11878),
            .in2(_gnd_net_),
            .in3(N__12348),
            .lcout(\spi_slave_1.bitcnt_rxe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_6_LC_4_2_0 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_6_LC_4_2_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_6_LC_4_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.num_leds_6_LC_4_2_0  (
            .in0(N__13693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.num_ledsZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27425),
            .ce(N__22362),
            .sr(N__27063));
    defparam \sb_translator_1.num_leds_5_LC_4_2_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_5_LC_4_2_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_5_LC_4_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_5_LC_4_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13855),
            .lcout(\sb_translator_1.num_ledsZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27425),
            .ce(N__22362),
            .sr(N__27063));
    defparam \sb_translator_1.num_leds_RNIN668_0_LC_4_3_0 .C_ON=1'b1;
    defparam \sb_translator_1.num_leds_RNIN668_0_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIN668_0_LC_4_3_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \sb_translator_1.num_leds_RNIN668_0_LC_4_3_0  (
            .in0(_gnd_net_),
            .in1(N__19104),
            .in2(N__19042),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.un1_num_leds_n_1 ),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_1_c_RNIDRFK_LC_4_3_1 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_1_c_RNIDRFK_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_1_c_RNIDRFK_LC_4_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_1_c_RNIDRFK_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__19041),
            .in2(N__19071),
            .in3(N__11023),
            .lcout(\sb_translator_1.un1_num_leds_n_2 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_1 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_2_c_RNIGVGK_LC_4_3_2 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_2_c_RNIGVGK_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_2_c_RNIGVGK_LC_4_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_2_c_RNIGVGK_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__19061),
            .in2(N__18685),
            .in3(N__11008),
            .lcout(\sb_translator_1.un1_num_leds_n_3 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_2 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_3_c_RNIJ3IK_LC_4_3_3 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_3_c_RNIJ3IK_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_3_c_RNIJ3IK_LC_4_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_3_c_RNIJ3IK_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__18680),
            .in2(N__18643),
            .in3(N__10996),
            .lcout(\sb_translator_1.un1_num_leds_n_4 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_3 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_4_c_RNIM7JK_LC_4_3_4 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_4_c_RNIM7JK_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_4_c_RNIM7JK_LC_4_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_4_c_RNIM7JK_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__18634),
            .in2(N__18402),
            .in3(N__10984),
            .lcout(\sb_translator_1.un1_num_leds_n_5 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_4 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_5_c_RNIPBKK_LC_4_3_5 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_5_c_RNIPBKK_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_5_c_RNIPBKK_LC_4_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_5_c_RNIPBKK_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__18392),
            .in2(N__18795),
            .in3(N__10969),
            .lcout(\sb_translator_1.un1_num_leds_n_6 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_5 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_6_c_RNISFLK_LC_4_3_6 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_6_c_RNISFLK_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_6_c_RNISFLK_LC_4_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_6_c_RNISFLK_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(N__18785),
            .in2(N__18753),
            .in3(N__10957),
            .lcout(\sb_translator_1.un1_num_leds_n_7 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_6 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_7_c_RNIVJMK_LC_4_3_7 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_7_c_RNIVJMK_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_7_c_RNIVJMK_LC_4_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_7_c_RNIVJMK_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__18749),
            .in2(N__18728),
            .in3(N__10942),
            .lcout(\sb_translator_1.un1_num_leds_n_8 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_7 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_8_c_RNI2ONK_LC_4_4_0 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_8_c_RNI2ONK_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_8_c_RNI2ONK_LC_4_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_8_c_RNI2ONK_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__18722),
            .in2(N__15934),
            .in3(N__11134),
            .lcout(\sb_translator_1.un1_num_leds_n_9 ),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_9_c_RNIC3RN_LC_4_4_1 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_9_c_RNIC3RN_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_9_c_RNIC3RN_LC_4_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_9_c_RNIC3RN_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__15932),
            .in2(N__15874),
            .in3(N__11122),
            .lcout(\sb_translator_1.un1_num_leds_n_10 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_9 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_10_c_RNITFLI_LC_4_4_2 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_10_c_RNITFLI_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_10_c_RNITFLI_LC_4_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_10_c_RNITFLI_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__15872),
            .in2(N__15901),
            .in3(N__11107),
            .lcout(\sb_translator_1.un1_num_leds_n_11 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_10 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_11_c_RNI0KMI_LC_4_4_3 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_11_c_RNI0KMI_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_11_c_RNI0KMI_LC_4_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_11_c_RNI0KMI_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__15900),
            .in2(N__20876),
            .in3(N__11095),
            .lcout(\sb_translator_1.un1_num_leds_n_12 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_11 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_12_c_RNI3ONI_LC_4_4_4 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_12_c_RNI3ONI_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_12_c_RNI3ONI_LC_4_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_12_c_RNI3ONI_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__20870),
            .in2(N__20775),
            .in3(N__11083),
            .lcout(\sb_translator_1.un1_num_leds_n_13 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_12 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_13_c_RNI6SOI_LC_4_4_5 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_13_c_RNI6SOI_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_13_c_RNI6SOI_LC_4_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_13_c_RNI6SOI_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__20765),
            .in2(N__20802),
            .in3(N__11071),
            .lcout(\sb_translator_1.un1_num_leds_n_14 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_13 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_14_c_RNI90QI_LC_4_4_6 .C_ON=1'b1;
    defparam \sb_translator_1.un1_num_leds_0_cry_14_c_RNI90QI_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_14_c_RNI90QI_LC_4_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_14_c_RNI90QI_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__20798),
            .in2(N__20962),
            .in3(N__11059),
            .lcout(\sb_translator_1.un1_num_leds_n_15 ),
            .ltout(),
            .carryin(\sb_translator_1.un1_num_leds_0_cry_14 ),
            .carryout(\sb_translator_1.un1_num_leds_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.un1_num_leds_0_cry_15_c_RNIQ9LB_LC_4_4_7 .C_ON=1'b0;
    defparam \sb_translator_1.un1_num_leds_0_cry_15_c_RNIQ9LB_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.un1_num_leds_0_cry_15_c_RNIQ9LB_LC_4_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \sb_translator_1.un1_num_leds_0_cry_15_c_RNIQ9LB_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__20961),
            .in2(_gnd_net_),
            .in3(N__11056),
            .lcout(\sb_translator_1.un1_num_leds_n_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.mosi_data_in_0_LC_4_5_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_0_LC_4_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_0_LC_4_5_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_0_LC_4_5_0  (
            .in0(N__11887),
            .in1(N__12228),
            .in2(_gnd_net_),
            .in3(N__12357),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_1_LC_4_5_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_1_LC_4_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_1_LC_4_5_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_1_LC_4_5_1  (
            .in0(N__12358),
            .in1(_gnd_net_),
            .in2(N__12244),
            .in3(N__13167),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_2_LC_4_5_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_2_LC_4_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_2_LC_4_5_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_2_LC_4_5_2  (
            .in0(N__11154),
            .in1(N__12232),
            .in2(_gnd_net_),
            .in3(N__12359),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_3_LC_4_5_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_3_LC_4_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_3_LC_4_5_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_3_LC_4_5_3  (
            .in0(N__12360),
            .in1(_gnd_net_),
            .in2(N__12245),
            .in3(N__12375),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_4_LC_4_5_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_4_LC_4_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_4_LC_4_5_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_4_LC_4_5_4  (
            .in0(N__12387),
            .in1(N__12236),
            .in2(_gnd_net_),
            .in3(N__12361),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_5_LC_4_5_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_5_LC_4_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_5_LC_4_5_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_5_LC_4_5_5  (
            .in0(N__12362),
            .in1(_gnd_net_),
            .in2(N__12246),
            .in3(N__13179),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_6_LC_4_5_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_6_LC_4_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_6_LC_4_5_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_6_LC_4_5_6  (
            .in0(N__13221),
            .in1(N__12240),
            .in2(_gnd_net_),
            .in3(N__12363),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \spi_slave_1.mosi_data_in_7_LC_4_5_7 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_7_LC_4_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_7_LC_4_5_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_7_LC_4_5_7  (
            .in0(N__12364),
            .in1(_gnd_net_),
            .in2(N__12247),
            .in3(N__13209),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27436),
            .ce(N__12063),
            .sr(N__27071));
    defparam \sb_translator_1.instr_tmp_5_LC_4_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_5_LC_4_6_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_5_LC_4_6_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \sb_translator_1.instr_tmp_5_LC_4_6_0  (
            .in0(N__22043),
            .in1(N__13848),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.instr_tmpZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27444),
            .ce(N__16971),
            .sr(N__27075));
    defparam \sb_translator_1.instr_tmp_6_LC_4_6_1 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_6_LC_4_6_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_6_LC_4_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sb_translator_1.instr_tmp_6_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__22042),
            .in2(_gnd_net_),
            .in3(N__13689),
            .lcout(\sb_translator_1.instr_tmpZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27444),
            .ce(N__16971),
            .sr(N__27075));
    defparam \sb_translator_1.instr_tmp_7_LC_4_6_2 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_7_LC_4_6_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_7_LC_4_6_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \sb_translator_1.instr_tmp_7_LC_4_6_2  (
            .in0(N__22044),
            .in1(N__13509),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.instr_tmpZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27444),
            .ce(N__16971),
            .sr(N__27075));
    defparam reset_n_input_RNIVGR4_LC_4_6_4.C_ON=1'b0;
    defparam reset_n_input_RNIVGR4_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam reset_n_input_RNIVGR4_LC_4_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_n_input_RNIVGR4_LC_4_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11281),
            .lcout(reset_n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_3_LC_4_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_3_LC_4_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_3_LC_4_7_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_we_3_LC_4_7_0  (
            .in0(N__13920),
            .in1(N__13947),
            .in2(N__17536),
            .in3(N__13301),
            .lcout(ram_we_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.ram_we_13_LC_4_7_1 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_13_LC_4_7_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_13_LC_4_7_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_we_13_LC_4_7_1  (
            .in0(N__17761),
            .in1(N__14048),
            .in2(N__11376),
            .in3(N__13919),
            .lcout(ram_we_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.cnt_RNILAHE_0_10_LC_4_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNILAHE_0_10_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNILAHE_0_10_LC_4_7_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \sb_translator_1.cnt_RNILAHE_0_10_LC_4_7_2  (
            .in0(N__17359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17311),
            .lcout(\sb_translator_1.cnt_RNILAHE_0Z0Z_10 ),
            .ltout(\sb_translator_1.cnt_RNILAHE_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_5_LC_4_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_5_LC_4_7_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_5_LC_4_7_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_we_5_LC_4_7_3  (
            .in0(N__13945),
            .in1(N__17794),
            .in2(N__11200),
            .in3(N__13921),
            .lcout(ram_we_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.ram_we_7_LC_4_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_7_LC_4_7_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_7_LC_4_7_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_we_7_LC_4_7_4  (
            .in0(N__13922),
            .in1(N__13946),
            .in2(N__17275),
            .in3(N__16950),
            .lcout(ram_we_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.ram_we_9_LC_4_7_5 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_9_LC_4_7_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_9_LC_4_7_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_we_9_LC_4_7_5  (
            .in0(N__16108),
            .in1(N__14283),
            .in2(N__11377),
            .in3(N__13923),
            .lcout(ram_we_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.cnt_RNILAHE_1_10_LC_4_7_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNILAHE_1_10_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNILAHE_1_10_LC_4_7_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \sb_translator_1.cnt_RNILAHE_1_10_LC_4_7_6  (
            .in0(N__17360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17312),
            .lcout(\sb_translator_1.cnt_RNILAHE_1Z0Z_10 ),
            .ltout(\sb_translator_1.cnt_RNILAHE_1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_11_LC_4_7_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_11_LC_4_7_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_11_LC_4_7_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_we_11_LC_4_7_7  (
            .in0(N__11369),
            .in1(N__16915),
            .in2(N__11356),
            .in3(N__13918),
            .lcout(ram_we_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27450),
            .ce(N__16785),
            .sr(N__27078));
    defparam \sb_translator_1.state_RNIHS98_0_LC_4_8_0 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIHS98_0_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIHS98_0_LC_4_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \sb_translator_1.state_RNIHS98_0_LC_4_8_0  (
            .in0(N__11329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22049),
            .lcout(\sb_translator_1.state_RNIHS98Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNIHS98_0_0_LC_4_8_1 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIHS98_0_0_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIHS98_0_0_LC_4_8_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \sb_translator_1.state_RNIHS98_0_0_LC_4_8_1  (
            .in0(N__22048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11328),
            .lcout(\sb_translator_1.state_RNIHS98_0Z0Z_0 ),
            .ltout(\sb_translator_1.state_RNIHS98_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_6_LC_4_8_2 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_6_LC_4_8_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_6_LC_4_8_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_sel_6_LC_4_8_2  (
            .in0(N__15841),
            .in1(N__21313),
            .in2(N__11338),
            .in3(N__16951),
            .lcout(ram_sel_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27457),
            .ce(N__17482),
            .sr(N__27083));
    defparam \sb_translator_1.state_RNIQIHP_0_LC_4_8_3 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIQIHP_0_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIQIHP_0_LC_4_8_3 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \sb_translator_1.state_RNIQIHP_0_LC_4_8_3  (
            .in0(N__22045),
            .in1(N__16860),
            .in2(_gnd_net_),
            .in3(N__22417),
            .lcout(\sb_translator_1.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNO_0_0_LC_4_8_4 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNO_0_0_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNO_0_0_LC_4_8_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \sb_translator_1.state_RNO_0_0_LC_4_8_4  (
            .in0(N__16862),
            .in1(N__22602),
            .in2(_gnd_net_),
            .in3(N__22046),
            .lcout(\sb_translator_1.N_729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNI9ILJ_0_LC_4_8_5 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNI9ILJ_0_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNI9ILJ_0_LC_4_8_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \sb_translator_1.state_RNI9ILJ_0_LC_4_8_5  (
            .in0(N__17232),
            .in1(N__22053),
            .in2(N__22603),
            .in3(N__11331),
            .lcout(\sb_translator_1.state_RNI9ILJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNI9ILJ_0_0_LC_4_8_6 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNI9ILJ_0_0_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNI9ILJ_0_0_LC_4_8_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \sb_translator_1.state_RNI9ILJ_0_0_LC_4_8_6  (
            .in0(N__11330),
            .in1(N__22598),
            .in2(N__22074),
            .in3(N__17233),
            .lcout(\sb_translator_1.state_RNI9ILJ_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNII30C_0_LC_4_8_7 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNII30C_0_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNII30C_0_LC_4_8_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \sb_translator_1.state_RNII30C_0_LC_4_8_7  (
            .in0(N__22047),
            .in1(_gnd_net_),
            .in2(N__17236),
            .in3(N__16861),
            .lcout(\sb_translator_1.state_RNII30CZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_a3_2_LC_4_9_0 .C_ON=1'b0;
    defparam \demux.N_418_i_0_a3_2_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_a3_2_LC_4_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \demux.N_418_i_0_a3_2_LC_4_9_0  (
            .in0(N__17947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11299),
            .lcout(),
            .ltout(\demux.N_877_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_9_LC_4_9_1 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_9_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_9_LC_4_9_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_418_i_0_o2_9_LC_4_9_1  (
            .in0(N__14485),
            .in1(N__11503),
            .in2(N__11494),
            .in3(N__11476),
            .lcout(\demux.N_418_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_6_LC_4_9_2 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_6_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_6_LC_4_9_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_418_i_0_o2_6_LC_4_9_2  (
            .in0(N__19645),
            .in1(N__11491),
            .in2(N__24360),
            .in3(N__11482),
            .lcout(\demux.N_418_i_0_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_a3_2_LC_4_9_3 .C_ON=1'b0;
    defparam \demux.N_421_i_0_a3_2_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_a3_2_LC_4_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_421_i_0_a3_2_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__11470),
            .in2(_gnd_net_),
            .in3(N__17946),
            .lcout(),
            .ltout(\demux.N_835_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_9_LC_4_9_4 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_9_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_9_LC_4_9_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_421_i_0_o2_9_LC_4_9_4  (
            .in0(N__11452),
            .in1(N__14484),
            .in2(N__11446),
            .in3(N__11425),
            .lcout(\demux.N_421_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_6_LC_4_9_5 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_6_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_6_LC_4_9_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_421_i_0_o2_6_LC_4_9_5  (
            .in0(N__11443),
            .in1(N__24349),
            .in2(N__11437),
            .in3(N__19643),
            .lcout(\demux.N_421_i_0_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_a3_1_LC_4_9_6 .C_ON=1'b0;
    defparam \demux.N_417_i_0_a3_1_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_a3_1_LC_4_9_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \demux.N_417_i_0_a3_1_LC_4_9_6  (
            .in0(N__19644),
            .in1(N__11419),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\demux.N_890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_a3_1_LC_4_9_7 .C_ON=1'b0;
    defparam \demux.N_423_i_0_a3_1_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_a3_1_LC_4_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_423_i_0_a3_1_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__11413),
            .in2(_gnd_net_),
            .in3(N__19642),
            .lcout(\demux.N_423_i_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_6_LC_4_10_0 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_6_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_6_LC_4_10_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_417_i_0_o2_6_LC_4_10_0  (
            .in0(N__17944),
            .in1(N__11407),
            .in2(N__21069),
            .in3(N__11389),
            .lcout(),
            .ltout(\demux.N_417_i_0_o2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_9_LC_4_10_1 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_9_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_9_LC_4_10_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_417_i_0_o2_9_LC_4_10_1  (
            .in0(N__11662),
            .in1(N__14471),
            .in2(N__11650),
            .in3(N__11647),
            .lcout(\demux.N_417_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_a3_1_LC_4_10_2 .C_ON=1'b0;
    defparam \demux.N_419_i_0_a3_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_a3_1_LC_4_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_419_i_0_a3_1_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__11641),
            .in2(_gnd_net_),
            .in3(N__19653),
            .lcout(\demux.N_419_i_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_6_LC_4_10_3 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_6_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_6_LC_4_10_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_419_i_0_o2_6_LC_4_10_3  (
            .in0(N__11635),
            .in1(N__17943),
            .in2(N__11623),
            .in3(N__21052),
            .lcout(),
            .ltout(\demux.N_419_i_0_o2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_9_LC_4_10_4 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_9_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_9_LC_4_10_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_419_i_0_o2_9_LC_4_10_4  (
            .in0(N__14470),
            .in1(N__11602),
            .in2(N__11587),
            .in3(N__11584),
            .lcout(\demux.N_419_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_a3_1_LC_4_10_5 .C_ON=1'b0;
    defparam \demux.N_420_i_0_a3_1_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_a3_1_LC_4_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \demux.N_420_i_0_a3_1_LC_4_10_5  (
            .in0(N__19654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11578),
            .lcout(\demux.N_420_i_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_6_LC_4_10_6 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_6_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_6_LC_4_10_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_420_i_0_o2_6_LC_4_10_6  (
            .in0(N__17945),
            .in1(N__11572),
            .in2(N__21070),
            .in3(N__11554),
            .lcout(),
            .ltout(\demux.N_420_i_0_o2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_9_LC_4_10_7 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_9_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_9_LC_4_10_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_420_i_0_o2_9_LC_4_10_7  (
            .in0(N__11542),
            .in1(N__14472),
            .in2(N__11533),
            .in3(N__11530),
            .lcout(\demux.N_420_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_6_LC_4_11_0 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_6_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_6_LC_4_11_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_slave_1.miso_data_out_6_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__23533),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.miso_data_outZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_1_LC_4_11_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_1_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_1_LC_4_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_1.miso_data_out_1_LC_4_11_1  (
            .in0(N__24022),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.miso_data_outZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_3_LC_4_11_2 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_3_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_3_LC_4_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_1.miso_data_out_3_LC_4_11_2  (
            .in0(N__24145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.miso_data_outZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_7_LC_4_11_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_7_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_7_LC_4_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_7_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23671),
            .lcout(\spi_slave_1.miso_data_outZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_18_LC_4_11_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_18_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_18_LC_4_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_18_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11749),
            .lcout(\spi_slave_1.miso_data_outZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_2_LC_4_11_6 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_2_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_2_LC_4_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_2_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17248),
            .lcout(\spi_slave_1.miso_data_outZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27481),
            .ce(N__14546),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_19_LC_4_12_0 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_19_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_19_LC_4_12_0 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \spi_slave_1.miso_RNO_19_LC_4_12_0  (
            .in0(N__11737),
            .in1(N__18571),
            .in2(N__11731),
            .in3(N__18521),
            .lcout(\spi_slave_1.m72_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_14_LC_4_12_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_14_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_14_LC_4_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_1.miso_data_out_14_LC_4_12_3  (
            .in0(N__14692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_1.miso_data_outZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27489),
            .ce(N__14539),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_13_LC_4_12_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_13_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_13_LC_4_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_13_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14698),
            .lcout(\spi_slave_1.miso_data_outZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27489),
            .ce(N__14539),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_12_LC_4_12_5 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_12_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_12_LC_4_12_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \spi_slave_1.miso_RNO_12_LC_4_12_5  (
            .in0(N__18522),
            .in1(N__11710),
            .in2(_gnd_net_),
            .in3(N__11704),
            .lcout(),
            .ltout(\spi_slave_1.miso_RNOZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_8_LC_4_12_6 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_8_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_8_LC_4_12_6 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \spi_slave_1.miso_RNO_8_LC_4_12_6  (
            .in0(N__11698),
            .in1(N__11943),
            .in2(N__11665),
            .in3(N__17962),
            .lcout(),
            .ltout(\spi_slave_1.m27_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_4_LC_4_12_7 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_4_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_4_LC_4_12_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \spi_slave_1.miso_RNO_4_LC_4_12_7  (
            .in0(N__11944),
            .in1(N__18604),
            .in2(N__11911),
            .in3(N__11908),
            .lcout(\spi_slave_1.N_28_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.mosi_buffer_1_LC_4_13_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_buffer_1_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_buffer_1_LC_4_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \spi_slave_1.mosi_buffer_1_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__11869),
            .in2(_gnd_net_),
            .in3(N__11776),
            .lcout(\spi_slave_1.mosi_bufferZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27494),
            .ce(),
            .sr(N__27114));
    defparam \spi_slave_1.mosi_buffer_0_LC_4_13_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_buffer_0_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_buffer_0_LC_4_13_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \spi_slave_1.mosi_buffer_0_LC_4_13_5  (
            .in0(N__11868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11791),
            .lcout(\spi_slave_1.mosi_bufferZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27494),
            .ce(),
            .sr(N__27114));
    defparam \spi_slave_1.mosi_data_in_10_LC_5_1_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_10_LC_5_1_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_10_LC_5_1_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_10_LC_5_1_0  (
            .in0(N__12045),
            .in1(N__12170),
            .in2(_gnd_net_),
            .in3(N__12349),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_11_LC_5_1_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_11_LC_5_1_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_11_LC_5_1_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_11_LC_5_1_1  (
            .in0(N__12350),
            .in1(_gnd_net_),
            .in2(N__12220),
            .in3(N__12003),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_12_LC_5_1_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_12_LC_5_1_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_12_LC_5_1_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_12_LC_5_1_2  (
            .in0(N__11991),
            .in1(N__12174),
            .in2(_gnd_net_),
            .in3(N__12351),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_13_LC_5_1_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_13_LC_5_1_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_13_LC_5_1_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_13_LC_5_1_3  (
            .in0(N__12352),
            .in1(_gnd_net_),
            .in2(N__12221),
            .in3(N__11979),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_14_LC_5_1_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_14_LC_5_1_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_14_LC_5_1_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_14_LC_5_1_4  (
            .in0(N__11967),
            .in1(N__12178),
            .in2(_gnd_net_),
            .in3(N__12353),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_15_LC_5_1_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_15_LC_5_1_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_15_LC_5_1_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_15_LC_5_1_5  (
            .in0(N__12354),
            .in1(_gnd_net_),
            .in2(N__12222),
            .in3(N__11955),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_16_LC_5_1_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_16_LC_5_1_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_16_LC_5_1_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_16_LC_5_1_6  (
            .in0(N__18438),
            .in1(N__12182),
            .in2(_gnd_net_),
            .in3(N__12355),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_in_17_LC_5_1_7 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_in_17_LC_5_1_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_in_17_LC_5_1_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \spi_slave_1.mosi_data_in_17_LC_5_1_7  (
            .in0(N__12356),
            .in1(_gnd_net_),
            .in2(N__12223),
            .in3(N__12399),
            .lcout(\spi_slave_1.mosi_data_inZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27426),
            .ce(N__12061),
            .sr(N__27064));
    defparam \spi_slave_1.mosi_data_out_9_LC_5_2_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_9_LC_5_2_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_9_LC_5_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_9_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12046),
            .lcout(mosi_data_out_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_8_LC_5_2_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_8_LC_5_2_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_8_LC_5_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_8_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12022),
            .lcout(mosi_data_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_10_LC_5_2_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_10_LC_5_2_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_10_LC_5_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_10_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12004),
            .lcout(mosi_data_out_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_11_LC_5_2_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_11_LC_5_2_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_11_LC_5_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_11_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11992),
            .lcout(mosi_data_out_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_12_LC_5_2_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_12_LC_5_2_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_12_LC_5_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_12_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11980),
            .lcout(mosi_data_out_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_13_LC_5_2_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_13_LC_5_2_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_13_LC_5_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_13_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11968),
            .lcout(mosi_data_out_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \spi_slave_1.mosi_data_out_14_LC_5_2_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_14_LC_5_2_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_14_LC_5_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_14_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11956),
            .lcout(mosi_data_out_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27428),
            .ce(N__18426),
            .sr(N__27066));
    defparam \sb_translator_1.num_leds_11_LC_5_3_0 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_11_LC_5_3_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_11_LC_5_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_11_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14644),
            .lcout(\sb_translator_1.num_ledsZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_12_LC_5_3_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_12_LC_5_3_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_12_LC_5_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_12_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22578),
            .lcout(\sb_translator_1.num_ledsZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_13_LC_5_3_2 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_13_LC_5_3_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_13_LC_5_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_13_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14605),
            .lcout(\sb_translator_1.num_ledsZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_14_LC_5_3_3 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_14_LC_5_3_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_14_LC_5_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_14_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22521),
            .lcout(\sb_translator_1.num_ledsZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_2_LC_5_3_4 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_2_LC_5_3_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_2_LC_5_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_2_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15961),
            .lcout(\sb_translator_1.num_ledsZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_3_LC_5_3_5 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_3_LC_5_3_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_3_LC_5_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_3_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17029),
            .lcout(\sb_translator_1.num_ledsZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_4_LC_5_3_6 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_4_LC_5_3_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_4_LC_5_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_4_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17002),
            .lcout(\sb_translator_1.num_ledsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_7_LC_5_3_7 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_7_LC_5_3_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_7_LC_5_3_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \sb_translator_1.num_leds_7_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__13513),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.num_ledsZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27432),
            .ce(N__22349),
            .sr(N__27068));
    defparam \sb_translator_1.num_leds_RNITOUT_8_LC_5_4_0 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNITOUT_8_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNITOUT_8_LC_5_4_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \sb_translator_1.num_leds_RNITOUT_8_LC_5_4_0  (
            .in0(N__20476),
            .in1(N__21356),
            .in2(N__15933),
            .in3(N__18717),
            .lcout(\sb_translator_1.num_leds_RNITOUTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNI0EVE_8_LC_5_4_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNI0EVE_8_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNI0EVE_8_LC_5_4_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \sb_translator_1.num_leds_RNI0EVE_8_LC_5_4_1  (
            .in0(N__18718),
            .in1(_gnd_net_),
            .in2(N__21364),
            .in3(N__15928),
            .lcout(\sb_translator_1.num_leds_RNI0EVEZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_8_LC_5_4_2 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_8_LC_5_4_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_8_LC_5_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.num_leds_8_LC_5_4_2  (
            .in0(N__12532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.num_ledsZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27437),
            .ce(N__22363),
            .sr(N__27072));
    defparam \sb_translator_1.num_leds_9_LC_5_4_3 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_9_LC_5_4_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_9_LC_5_4_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \sb_translator_1.num_leds_9_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__12484),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.num_ledsZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27437),
            .ce(N__22363),
            .sr(N__27072));
    defparam \sb_translator_1.addr_out_RNO_0_0_LC_5_4_4 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_0_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_0_LC_5_4_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_0_LC_5_4_4  (
            .in0(N__12531),
            .in1(N__22997),
            .in2(_gnd_net_),
            .in3(N__12517),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_RNO_0_1_LC_5_4_5 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_1_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_1_LC_5_4_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_1_LC_5_4_5  (
            .in0(N__22998),
            .in1(N__12483),
            .in2(_gnd_net_),
            .in3(N__12472),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_RNO_0_2_LC_5_4_6 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_2_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_2_LC_5_4_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_2_LC_5_4_6  (
            .in0(N__12414),
            .in1(N__22999),
            .in2(_gnd_net_),
            .in3(N__12442),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_10_LC_5_4_7 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_10_LC_5_4_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_10_LC_5_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_10_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12415),
            .lcout(\sb_translator_1.num_ledsZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27437),
            .ce(N__22363),
            .sr(N__27072));
    defparam \spi_slave_1.mosi_data_out_16_LC_5_5_0 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_16_LC_5_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_16_LC_5_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_16_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12403),
            .lcout(mosi_data_out_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_3_LC_5_5_1 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_3_LC_5_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_3_LC_5_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_3_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12388),
            .lcout(mosi_data_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_2_LC_5_5_2 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_2_LC_5_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_2_LC_5_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_2_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12376),
            .lcout(mosi_data_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_5_LC_5_5_3 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_5_LC_5_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_5_LC_5_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_5_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13222),
            .lcout(mosi_data_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_6_LC_5_5_4 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_6_LC_5_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_6_LC_5_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_6_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13210),
            .lcout(mosi_data_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_7_LC_5_5_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_7_LC_5_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_7_LC_5_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_7_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13194),
            .lcout(mosi_data_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_4_LC_5_5_6 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_4_LC_5_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_4_LC_5_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_4_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13180),
            .lcout(mosi_data_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \spi_slave_1.mosi_data_out_0_LC_5_5_7 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_0_LC_5_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_0_LC_5_5_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_slave_1.mosi_data_out_0_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__13168),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(mosi_data_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27445),
            .ce(N__18425),
            .sr(N__27076));
    defparam \sb_translator_1.data_out_0_LC_5_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_0_LC_5_6_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_0_LC_5_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sb_translator_1.data_out_0_LC_5_6_0  (
            .in0(N__16022),
            .in1(N__21993),
            .in2(_gnd_net_),
            .in3(N__16003),
            .lcout(ram_data_in_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_1_LC_5_6_1 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_1_LC_5_6_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_1_LC_5_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.data_out_1_LC_5_6_1  (
            .in0(N__21989),
            .in1(N__15967),
            .in2(_gnd_net_),
            .in3(N__15989),
            .lcout(ram_data_in_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_2_LC_5_6_2 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_2_LC_5_6_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_2_LC_5_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \sb_translator_1.data_out_2_LC_5_6_2  (
            .in0(N__15940),
            .in1(N__15956),
            .in2(_gnd_net_),
            .in3(N__21994),
            .lcout(ram_data_in_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_3_LC_5_6_3 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_3_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_3_LC_5_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.data_out_3_LC_5_6_3  (
            .in0(N__21990),
            .in1(N__17008),
            .in2(_gnd_net_),
            .in3(N__17024),
            .lcout(ram_data_in_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_4_LC_5_6_4 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_4_LC_5_6_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_4_LC_5_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sb_translator_1.data_out_4_LC_5_6_4  (
            .in0(N__17000),
            .in1(N__21995),
            .in2(_gnd_net_),
            .in3(N__16981),
            .lcout(ram_data_in_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_5_LC_5_6_5 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_5_LC_5_6_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_5_LC_5_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.data_out_5_LC_5_6_5  (
            .in0(N__21991),
            .in1(N__13861),
            .in2(_gnd_net_),
            .in3(N__13847),
            .lcout(ram_data_in_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_6_LC_5_6_6 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_6_LC_5_6_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_6_LC_5_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \sb_translator_1.data_out_6_LC_5_6_6  (
            .in0(N__13702),
            .in1(N__13688),
            .in2(_gnd_net_),
            .in3(N__21996),
            .lcout(ram_data_in_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.data_out_7_LC_5_6_7 .C_ON=1'b0;
    defparam \sb_translator_1.data_out_7_LC_5_6_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.data_out_7_LC_5_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.data_out_7_LC_5_6_7  (
            .in0(N__21992),
            .in1(N__13519),
            .in2(_gnd_net_),
            .in3(N__13508),
            .lcout(ram_data_in_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27451),
            .ce(N__16789),
            .sr(N__27079));
    defparam \sb_translator_1.ram_we_0_LC_5_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_0_LC_5_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_0_LC_5_7_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_we_0_LC_5_7_0  (
            .in0(N__14011),
            .in1(N__16099),
            .in2(N__17728),
            .in3(N__13990),
            .lcout(ram_we_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_2_LC_5_7_1 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_2_LC_5_7_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_2_LC_5_7_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_we_2_LC_5_7_1  (
            .in0(N__13987),
            .in1(N__17529),
            .in2(N__13306),
            .in3(N__14014),
            .lcout(ram_we_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_10_LC_5_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_10_LC_5_7_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_10_LC_5_7_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_we_10_LC_5_7_2  (
            .in0(N__13250),
            .in1(N__13302),
            .in2(N__16918),
            .in3(N__13991),
            .lcout(ram_we_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_8_LC_5_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_8_LC_5_7_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_8_LC_5_7_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_we_8_LC_5_7_3  (
            .in0(N__13989),
            .in1(N__13254),
            .in2(N__16104),
            .in3(N__14282),
            .lcout(ram_we_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_12_LC_5_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_12_LC_5_7_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_12_LC_5_7_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_we_12_LC_5_7_4  (
            .in0(N__17757),
            .in1(N__14049),
            .in2(N__13255),
            .in3(N__13992),
            .lcout(ram_we_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_4_LC_5_7_5 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_4_LC_5_7_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_4_LC_5_7_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_we_4_LC_5_7_5  (
            .in0(N__13988),
            .in1(N__17792),
            .in2(N__14053),
            .in3(N__14012),
            .lcout(ram_we_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_6_LC_5_7_6 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_6_LC_5_7_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_6_LC_5_7_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_we_6_LC_5_7_6  (
            .in0(N__14013),
            .in1(N__16945),
            .in2(N__17265),
            .in3(N__13993),
            .lcout(ram_we_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_we_1_LC_5_7_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_1_LC_5_7_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_we_1_LC_5_7_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_we_1_LC_5_7_7  (
            .in0(N__17727),
            .in1(N__13951),
            .in2(N__16103),
            .in3(N__13924),
            .lcout(ram_we_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27458),
            .ce(N__16784),
            .sr(N__27084));
    defparam \sb_translator_1.ram_sel_11_LC_5_8_0 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_11_LC_5_8_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_11_LC_5_8_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_11_LC_5_8_0  (
            .in0(N__16071),
            .in1(N__16916),
            .in2(N__13873),
            .in3(N__14343),
            .lcout(ram_sel_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27466),
            .ce(N__17483),
            .sr(N__27089));
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_9_LC_5_8_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_9_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_9_LC_5_8_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \sb_translator_1.cnt_leds_RNI1VFQ_9_LC_5_8_1  (
            .in0(N__21362),
            .in1(_gnd_net_),
            .in2(N__21418),
            .in3(N__22052),
            .lcout(\sb_translator_1.N_1091 ),
            .ltout(\sb_translator_1.N_1091_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_13_LC_5_8_2 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_13_LC_5_8_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_13_LC_5_8_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_sel_13_LC_5_8_2  (
            .in0(N__17750),
            .in1(N__15809),
            .in2(N__13879),
            .in3(N__14344),
            .lcout(ram_sel_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27466),
            .ce(N__17483),
            .sr(N__27089));
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_0_9_LC_5_8_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_0_9_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_0_9_LC_5_8_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \sb_translator_1.cnt_leds_RNI1VFQ_0_9_LC_5_8_3  (
            .in0(N__21361),
            .in1(_gnd_net_),
            .in2(N__21417),
            .in3(N__22051),
            .lcout(\sb_translator_1.N_1089 ),
            .ltout(\sb_translator_1.N_1089_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_10_LC_5_8_4 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_10_LC_5_8_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_10_LC_5_8_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_10_LC_5_8_4  (
            .in0(N__16070),
            .in1(N__14295),
            .in2(N__13876),
            .in3(N__16917),
            .lcout(ram_sel_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27466),
            .ce(N__17483),
            .sr(N__27089));
    defparam \sb_translator_1.ram_sel_9_LC_5_8_5 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_9_LC_5_8_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_9_LC_5_8_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_9_LC_5_8_5  (
            .in0(N__14342),
            .in1(N__16038),
            .in2(N__14281),
            .in3(N__13872),
            .lcout(ram_sel_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27466),
            .ce(N__17483),
            .sr(N__27089));
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_1_9_LC_5_8_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_1_9_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_1_9_LC_5_8_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \sb_translator_1.cnt_leds_RNI1VFQ_1_9_LC_5_8_6  (
            .in0(N__22050),
            .in1(N__21409),
            .in2(_gnd_net_),
            .in3(N__21360),
            .lcout(\sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9 ),
            .ltout(\sb_translator_1.cnt_leds_RNI1VFQ_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_7_LC_5_8_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_7_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_7_LC_5_8_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \sb_translator_1.ram_sel_7_LC_5_8_7  (
            .in0(N__14341),
            .in1(N__16946),
            .in2(N__14218),
            .in3(N__15840),
            .lcout(ram_sel_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27466),
            .ce(N__17483),
            .sr(N__27089));
    defparam \demux.N_422_i_0_o2_6_LC_5_9_0 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_6_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_6_LC_5_9_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_422_i_0_o2_6_LC_5_9_0  (
            .in0(N__14215),
            .in1(N__21060),
            .in2(N__14200),
            .in3(N__17936),
            .lcout(),
            .ltout(\demux.N_422_i_0_o2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_9_LC_5_9_1 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_9_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_9_LC_5_9_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_422_i_0_o2_9_LC_5_9_1  (
            .in0(N__14182),
            .in1(N__14477),
            .in2(N__14170),
            .in3(N__14104),
            .lcout(\demux.N_422_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_6_LC_5_9_2 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_6_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_6_LC_5_9_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_423_i_0_o2_6_LC_5_9_2  (
            .in0(N__14167),
            .in1(N__21059),
            .in2(N__14152),
            .in3(N__17935),
            .lcout(),
            .ltout(\demux.N_423_i_0_o2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_9_LC_5_9_3 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_9_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_9_LC_5_9_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_423_i_0_o2_9_LC_5_9_3  (
            .in0(N__14137),
            .in1(N__14476),
            .in2(N__14125),
            .in3(N__14122),
            .lcout(\demux.N_423_i_0_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_a3_1_LC_5_9_4 .C_ON=1'b0;
    defparam \demux.N_422_i_0_a3_1_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_a3_1_LC_5_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_422_i_0_a3_1_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__14116),
            .in2(_gnd_net_),
            .in3(N__19651),
            .lcout(\demux.N_422_i_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_6_0_LC_5_9_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_6_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_6_0_LC_5_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_424_i_0_o2_6_0_LC_5_9_5  (
            .in0(N__17937),
            .in1(N__14098),
            .in2(N__21071),
            .in3(N__14083),
            .lcout(),
            .ltout(\demux.N_424_i_0_o2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_9_0_LC_5_9_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_9_0_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_9_0_LC_5_9_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_424_i_0_o2_9_0_LC_5_9_6  (
            .in0(N__14478),
            .in1(N__14071),
            .in2(N__14056),
            .in3(N__14371),
            .lcout(\demux.N_424_i_0_o2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a3_1_LC_5_9_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a3_1_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a3_1_LC_5_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \demux.N_424_i_0_a3_1_LC_5_9_7  (
            .in0(N__19652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14383),
            .lcout(\demux.N_424_i_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_0_LC_5_10_0 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_0_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_0_LC_5_10_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_0_LC_5_10_0  (
            .in0(N__21310),
            .in1(N__17719),
            .in2(N__16054),
            .in3(N__14310),
            .lcout(ram_sel_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_2_LC_5_10_1 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_2_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_2_LC_5_10_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_2_LC_5_10_1  (
            .in0(N__14312),
            .in1(N__21312),
            .in2(N__17527),
            .in3(N__16077),
            .lcout(ram_sel_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_1_LC_5_10_2 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_1_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_1_LC_5_10_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_1_LC_5_10_2  (
            .in0(N__14364),
            .in1(N__14346),
            .in2(N__16053),
            .in3(N__17720),
            .lcout(ram_sel_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_3_LC_5_10_3 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_3_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_3_LC_5_10_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_3_LC_5_10_3  (
            .in0(N__14345),
            .in1(N__14365),
            .in2(N__17528),
            .in3(N__16078),
            .lcout(ram_sel_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_5_LC_5_10_4 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_5_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_5_LC_5_10_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_sel_5_LC_5_10_4  (
            .in0(N__14363),
            .in1(N__17788),
            .in2(N__14350),
            .in3(N__15819),
            .lcout(ram_sel_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_4_LC_5_10_5 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_4_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_4_LC_5_10_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_4_LC_5_10_5  (
            .in0(N__14313),
            .in1(N__21311),
            .in2(N__17793),
            .in3(N__15820),
            .lcout(ram_sel_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_12_LC_5_10_6 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_12_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_12_LC_5_10_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \sb_translator_1.ram_sel_12_LC_5_10_6  (
            .in0(N__17749),
            .in1(N__15818),
            .in2(N__14233),
            .in3(N__14311),
            .lcout(ram_sel_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \sb_translator_1.ram_sel_8_LC_5_10_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_8_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.ram_sel_8_LC_5_10_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \sb_translator_1.ram_sel_8_LC_5_10_7  (
            .in0(N__14314),
            .in1(N__16049),
            .in2(N__14284),
            .in3(N__14232),
            .lcout(ram_sel_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27482),
            .ce(N__17494),
            .sr(N__27101));
    defparam \demux.N_424_i_0_o2_11_LC_5_11_0 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_11_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_11_LC_5_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \demux.N_424_i_0_o2_11_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__17854),
            .in2(_gnd_net_),
            .in3(N__17875),
            .lcout(\demux.N_236 ),
            .ltout(\demux.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_16_LC_5_11_1 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_16_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_16_LC_5_11_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \demux.N_424_i_0_o2_16_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__14436),
            .in2(N__14491),
            .in3(N__14415),
            .lcout(\demux.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_14_LC_5_11_2 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_14_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_14_LC_5_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \demux.N_424_i_0_o2_14_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__19806),
            .in2(_gnd_net_),
            .in3(N__19752),
            .lcout(\demux.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_10_LC_5_11_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_10_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_10_LC_5_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \demux.N_424_i_0_o2_10_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__14437),
            .in2(_gnd_net_),
            .in3(N__14416),
            .lcout(\demux.N_235 ),
            .ltout(\demux.N_235_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_2_LC_5_11_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_2_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_2_LC_5_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \demux.N_424_i_0_a2_2_LC_5_11_4  (
            .in0(N__17857),
            .in1(N__17879),
            .in2(N__14488),
            .in3(N__17891),
            .lcout(\demux.N_424_i_0_a2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_6_LC_5_11_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_6_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_6_LC_5_11_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \demux.N_424_i_0_a2_6_LC_5_11_5  (
            .in0(N__17893),
            .in1(N__14442),
            .in2(N__19602),
            .in3(N__14419),
            .lcout(\demux.N_424_i_0_a2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_0_LC_5_11_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_0_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_0_LC_5_11_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \demux.N_424_i_0_a2_0_LC_5_11_6  (
            .in0(N__14418),
            .in1(N__19595),
            .in2(N__14443),
            .in3(N__17892),
            .lcout(\demux.N_424_i_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_2_LC_5_11_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_2_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_2_LC_5_11_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \demux.N_424_i_0_o2_0_2_LC_5_11_7  (
            .in0(N__17855),
            .in1(N__14438),
            .in2(N__17881),
            .in3(N__14417),
            .lcout(\demux.N_424_i_0_o2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_0_LC_5_12_0 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_0_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_0_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17806),
            .lcout(\spi_slave_1.miso_data_outZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_9_LC_5_12_1 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_9_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_9_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_9_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14398),
            .lcout(\spi_slave_1.miso_data_outZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_10_LC_5_12_2 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_10_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_10_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_10_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14509),
            .lcout(\spi_slave_1.miso_data_outZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_11_LC_5_12_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_11_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_11_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_11_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14503),
            .lcout(\spi_slave_1.miso_data_outZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_12_LC_5_12_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_12_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_12_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_12_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14497),
            .lcout(\spi_slave_1.miso_data_outZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_15_LC_5_12_5 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_15_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_15_LC_5_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_15_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14686),
            .lcout(\spi_slave_1.miso_data_outZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_16_LC_5_12_6 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_16_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_16_LC_5_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_16_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14680),
            .lcout(\spi_slave_1.miso_data_outZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_data_out_17_LC_5_12_7 .C_ON=1'b0;
    defparam \spi_slave_1.miso_data_out_17_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \spi_slave_1.miso_data_out_17_LC_5_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.miso_data_out_17_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14650),
            .lcout(\spi_slave_1.miso_data_outZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27495),
            .ce(N__14551),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_out_10_LC_5_13_0 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_10_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_10_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_10_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15189),
            .lcout(miso_data_in_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_11_LC_5_13_1 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_11_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_11_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_11_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14973),
            .lcout(miso_data_in_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_12_LC_5_13_2 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_12_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_12_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_12_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14769),
            .lcout(miso_data_in_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_13_LC_5_13_3 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_13_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_13_LC_5_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_13_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16590),
            .lcout(miso_data_in_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_14_LC_5_13_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_14_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_14_LC_5_13_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \sb_translator_1.instr_out_14_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__16386),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(miso_data_in_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_15_LC_5_13_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_15_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_15_LC_5_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_15_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16170),
            .lcout(miso_data_in_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_16_LC_5_13_6 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_16_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_16_LC_5_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_16_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18057),
            .lcout(miso_data_in_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.instr_out_17_LC_5_13_7 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_17_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_17_LC_5_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.instr_out_17_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14674),
            .lcout(miso_data_in_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27499),
            .ce(N__23994),
            .sr(N__27124));
    defparam \sb_translator_1.addr_out_RNO_0_3_LC_6_2_0 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_3_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_3_LC_6_2_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_3_LC_6_2_0  (
            .in0(N__14643),
            .in1(N__23009),
            .in2(_gnd_net_),
            .in3(N__14632),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_RNO_0_5_LC_6_2_1 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_5_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_5_LC_6_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_5_LC_6_2_1  (
            .in0(N__23010),
            .in1(N__14604),
            .in2(_gnd_net_),
            .in3(N__14593),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_0_LC_6_3_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_0_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_0_LC_6_3_0 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \sb_translator_1.cnt_leds_RNIO2NL_0_0_LC_6_3_0  (
            .in0(N__19095),
            .in1(N__18966),
            .in2(N__19037),
            .in3(N__18994),
            .lcout(\sb_translator_1.state56_a_5_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_0_LC_6_3_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_0_LC_6_3_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_0_LC_6_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_0_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16024),
            .lcout(\sb_translator_1.cnt19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27438),
            .ce(N__22348),
            .sr(N__27073));
    defparam \sb_translator_1.num_leds_1_LC_6_3_2 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_1_LC_6_3_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_1_LC_6_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_1_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15997),
            .lcout(\sb_translator_1.num_ledsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27438),
            .ce(N__22348),
            .sr(N__27073));
    defparam \sb_translator_1.cnt_ram_read_RNIPFJ32_1_LC_6_3_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNIPFJ32_1_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNIPFJ32_1_LC_6_3_3 .LUT_INIT=16'b1111111100010101;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNIPFJ32_1_LC_6_3_3  (
            .in0(N__22405),
            .in1(N__17451),
            .in2(N__17418),
            .in3(N__22259),
            .lcout(\sb_translator_1.cnt_ram_read_RNIPFJ32Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_0_1_LC_6_3_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_0_1_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_0_1_LC_6_3_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNINT0G1_0_1_LC_6_3_4  (
            .in0(N__17447),
            .in1(N__17402),
            .in2(_gnd_net_),
            .in3(N__22401),
            .lcout(\sb_translator_1.send_leds_n_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_LC_6_3_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_LC_6_3_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNINT0G1_1_LC_6_3_5  (
            .in0(N__22403),
            .in1(_gnd_net_),
            .in2(N__17417),
            .in3(N__17450),
            .lcout(\sb_translator_1.cnt_ram_read_RNINT0G1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_1_LC_6_3_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_1_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_1_1_LC_6_3_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNINT0G1_1_1_LC_6_3_6  (
            .in0(N__17448),
            .in1(N__17406),
            .in2(_gnd_net_),
            .in3(N__22402),
            .lcout(\sb_translator_1.cnt_ram_read_RNINT0G1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_2_1_LC_6_3_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_2_1_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNINT0G1_2_1_LC_6_3_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNINT0G1_2_1_LC_6_3_7  (
            .in0(N__22404),
            .in1(_gnd_net_),
            .in2(N__17416),
            .in3(N__17449),
            .lcout(\sb_translator_1.cnt_ram_read_RNINT0G1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIH2E91_9_LC_6_4_0 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIH2E91_9_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIH2E91_9_LC_6_4_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \sb_translator_1.num_leds_RNIH2E91_9_LC_6_4_0  (
            .in0(N__20436),
            .in1(N__15923),
            .in2(N__15873),
            .in3(N__19181),
            .lcout(\sb_translator_1.num_leds_RNIH2E91Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIRUGT_10_LC_6_4_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIRUGT_10_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIRUGT_10_LC_6_4_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \sb_translator_1.num_leds_RNIRUGT_10_LC_6_4_1  (
            .in0(N__15895),
            .in1(N__15868),
            .in2(_gnd_net_),
            .in3(N__19148),
            .lcout(\sb_translator_1.num_leds_RNIRUGTZ0Z_10 ),
            .ltout(\sb_translator_1.num_leds_RNIRUGTZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIP02R1_11_LC_6_4_2 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIP02R1_11_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIP02R1_11_LC_6_4_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.num_leds_RNIP02R1_11_LC_6_4_2  (
            .in0(N__20865),
            .in1(N__21387),
            .in2(N__14701),
            .in3(N__15894),
            .lcout(\sb_translator_1.num_leds_RNIP02R1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIU1HT_11_LC_6_4_3 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIU1HT_11_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIU1HT_11_LC_6_4_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \sb_translator_1.num_leds_RNIU1HT_11_LC_6_4_3  (
            .in0(N__15896),
            .in1(_gnd_net_),
            .in2(N__21398),
            .in3(N__20866),
            .lcout(\sb_translator_1.num_leds_RNIU1HTZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIHKEQ_9_LC_6_4_4 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIHKEQ_9_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIHKEQ_9_LC_6_4_4 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \sb_translator_1.num_leds_RNIHKEQ_9_LC_6_4_4  (
            .in0(N__15867),
            .in1(N__15924),
            .in2(_gnd_net_),
            .in3(N__19180),
            .lcout(\sb_translator_1.num_leds_RNIHKEQZ0Z_9 ),
            .ltout(\sb_translator_1.num_leds_RNIHKEQZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNICJVN1_10_LC_6_4_5 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNICJVN1_10_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNICJVN1_10_LC_6_4_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.num_leds_RNICJVN1_10_LC_6_4_5  (
            .in0(N__15893),
            .in1(N__15863),
            .in2(N__15844),
            .in3(N__19147),
            .lcout(\sb_translator_1.num_leds_RNICJVN1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI39BU_10_LC_6_4_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI39BU_10_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI39BU_10_LC_6_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \sb_translator_1.cnt_leds_RNI39BU_10_LC_6_4_6  (
            .in0(N__19150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19183),
            .lcout(\sb_translator_1.ram_sel_6_0_0_a2_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI39BU_0_10_LC_6_4_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI39BU_0_10_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI39BU_0_10_LC_6_4_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \sb_translator_1.cnt_leds_RNI39BU_0_10_LC_6_4_7  (
            .in0(N__19182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19149),
            .lcout(\sb_translator_1.cnt_leds_RNI39BU_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_0_LC_6_5_0 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_0_LC_6_5_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_0_LC_6_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_0_LC_6_5_0  (
            .in0(N__15790),
            .in1(N__22203),
            .in2(_gnd_net_),
            .in3(N__18997),
            .lcout(addr_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_1_LC_6_5_1 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_1_LC_6_5_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_1_LC_6_5_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \sb_translator_1.addr_out_1_LC_6_5_1  (
            .in0(N__22199),
            .in1(_gnd_net_),
            .in2(N__15571),
            .in3(N__18970),
            .lcout(addr_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_2_LC_6_5_2 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_2_LC_6_5_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_2_LC_6_5_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \sb_translator_1.addr_out_2_LC_6_5_2  (
            .in0(N__18940),
            .in1(N__22204),
            .in2(_gnd_net_),
            .in3(N__15355),
            .lcout(addr_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_3_LC_6_5_3 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_3_LC_6_5_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_3_LC_6_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_3_LC_6_5_3  (
            .in0(N__22200),
            .in1(N__15139),
            .in2(_gnd_net_),
            .in3(N__18915),
            .lcout(addr_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_4_LC_6_5_4 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_4_LC_6_5_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_4_LC_6_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_4_LC_6_5_4  (
            .in0(N__22537),
            .in1(N__22205),
            .in2(_gnd_net_),
            .in3(N__18888),
            .lcout(addr_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_5_LC_6_5_5 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_5_LC_6_5_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_5_LC_6_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_5_LC_6_5_5  (
            .in0(N__22201),
            .in1(N__16759),
            .in2(_gnd_net_),
            .in3(N__18857),
            .lcout(addr_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_6_LC_6_5_6 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_6_LC_6_5_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_6_LC_6_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_6_LC_6_5_6  (
            .in0(N__22483),
            .in1(N__22206),
            .in2(_gnd_net_),
            .in3(N__18830),
            .lcout(addr_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.addr_out_7_LC_6_5_7 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_7_LC_6_5_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_7_LC_6_5_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \sb_translator_1.addr_out_7_LC_6_5_7  (
            .in0(N__22202),
            .in1(_gnd_net_),
            .in2(N__22900),
            .in3(N__19244),
            .lcout(addr_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27452),
            .ce(N__18027),
            .sr(N__27080));
    defparam \sb_translator_1.cnt_RNILAHE_2_10_LC_6_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNILAHE_2_10_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNILAHE_2_10_LC_6_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \sb_translator_1.cnt_RNILAHE_2_10_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__17367),
            .in2(_gnd_net_),
            .in3(N__17319),
            .lcout(\sb_translator_1.cnt_RNILAHE_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI39BU_1_10_LC_6_6_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI39BU_1_10_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI39BU_1_10_LC_6_6_1 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \sb_translator_1.cnt_leds_RNI39BU_1_10_LC_6_6_1  (
            .in0(N__19185),
            .in1(N__19152),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_leds_RNI39BU_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI39BU_2_10_LC_6_6_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI39BU_2_10_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI39BU_2_10_LC_6_6_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \sb_translator_1.cnt_leds_RNI39BU_2_10_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__19184),
            .in2(_gnd_net_),
            .in3(N__19153),
            .lcout(\sb_translator_1.cnt_leds_RNI39BU_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_tmp_0_LC_6_6_3 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_0_LC_6_6_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_0_LC_6_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sb_translator_1.instr_tmp_0_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__16023),
            .in2(_gnd_net_),
            .in3(N__22015),
            .lcout(\sb_translator_1.instr_tmpZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27459),
            .ce(N__16975),
            .sr(N__27085));
    defparam \sb_translator_1.instr_tmp_1_LC_6_6_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_1_LC_6_6_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_1_LC_6_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \sb_translator_1.instr_tmp_1_LC_6_6_4  (
            .in0(N__22013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15996),
            .lcout(\sb_translator_1.instr_tmpZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27459),
            .ce(N__16975),
            .sr(N__27085));
    defparam \sb_translator_1.instr_tmp_2_LC_6_6_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_2_LC_6_6_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_2_LC_6_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sb_translator_1.instr_tmp_2_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__15957),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(\sb_translator_1.instr_tmpZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27459),
            .ce(N__16975),
            .sr(N__27085));
    defparam \sb_translator_1.instr_tmp_3_LC_6_6_6 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_3_LC_6_6_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_3_LC_6_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \sb_translator_1.instr_tmp_3_LC_6_6_6  (
            .in0(N__22014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17025),
            .lcout(\sb_translator_1.instr_tmpZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27459),
            .ce(N__16975),
            .sr(N__27085));
    defparam \sb_translator_1.instr_tmp_4_LC_6_6_7 .C_ON=1'b0;
    defparam \sb_translator_1.instr_tmp_4_LC_6_6_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_tmp_4_LC_6_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sb_translator_1.instr_tmp_4_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__17001),
            .in2(_gnd_net_),
            .in3(N__22017),
            .lcout(\sb_translator_1.instr_tmpZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27459),
            .ce(N__16975),
            .sr(N__27085));
    defparam \sb_translator_1.rgb_data_tmp_18_LC_6_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_18_LC_6_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_18_LC_6_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_18_LC_6_7_0  (
            .in0(N__20994),
            .in1(N__21615),
            .in2(N__21576),
            .in3(N__21541),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27467),
            .ce(N__25058),
            .sr(N__27090));
    defparam \sb_translator_1.rgb_data_tmp_16_LC_6_7_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_16_LC_6_7_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_16_LC_6_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_16_LC_6_7_1  (
            .in0(N__20002),
            .in1(N__19940),
            .in2(N__19970),
            .in3(N__19895),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27467),
            .ce(N__25058),
            .sr(N__27090));
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_7_LC_6_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_7_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_7_LC_6_7_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \sb_translator_1.ram_we_6_0_0_a2_1_7_LC_6_7_2  (
            .in0(N__17629),
            .in1(N__17576),
            .in2(_gnd_net_),
            .in3(N__17681),
            .lcout(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_6_0_0_a2_2_11_LC_6_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_6_0_0_a2_2_11_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_we_6_0_0_a2_2_11_LC_6_7_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \sb_translator_1.ram_we_6_0_0_a2_2_11_LC_6_7_3  (
            .in0(N__17682),
            .in1(N__17630),
            .in2(_gnd_net_),
            .in3(N__17577),
            .lcout(\sb_translator_1.ram_we_6_0_0_a2_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNIEL0N9_0_6_LC_6_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIEL0N9_0_6_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIEL0N9_0_6_LC_6_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.state_RNIEL0N9_0_6_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16888),
            .lcout(\sb_translator_1.state_RNIEL0N9_0Z0Z_6 ),
            .ltout(\sb_translator_1.state_RNIEL0N9_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNIOH7V9_0_LC_6_7_5 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNIOH7V9_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNIOH7V9_0_LC_6_7_5 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \sb_translator_1.state_RNIOH7V9_0_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__22009),
            .in2(N__16867),
            .in3(N__16863),
            .lcout(\sb_translator_1.state_RNIOH7V9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNI88IGA_0_LC_6_7_7 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNI88IGA_0_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNI88IGA_0_LC_6_7_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \sb_translator_1.state_RNI88IGA_0_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(N__17493),
            .in2(_gnd_net_),
            .in3(N__17458),
            .lcout(\sb_translator_1.state_RNI88IGAZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_0_LC_6_8_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_0_LC_6_8_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_ram_read_0_LC_6_8_0 .LUT_INIT=16'b0000000001000001;
    LogicCell40 \sb_translator_1.cnt_ram_read_0_LC_6_8_0  (
            .in0(N__27208),
            .in1(N__22421),
            .in2(N__17452),
            .in3(N__22306),
            .lcout(\sb_translator_1.cnt_ram_readZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27474),
            .ce(),
            .sr(N__27096));
    defparam \sb_translator_1.cnt_ram_read_1_LC_6_8_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_1_LC_6_8_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_ram_read_1_LC_6_8_1 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \sb_translator_1.cnt_ram_read_1_LC_6_8_1  (
            .in0(N__22422),
            .in1(N__17443),
            .in2(N__17419),
            .in3(N__17812),
            .lcout(\sb_translator_1.cnt_ram_readZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27474),
            .ce(),
            .sr(N__27096));
    defparam \sb_translator_1.state_leds_LC_6_8_2 .C_ON=1'b0;
    defparam \sb_translator_1.state_leds_LC_6_8_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.state_leds_LC_6_8_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \sb_translator_1.state_leds_LC_6_8_2  (
            .in0(N__27207),
            .in1(N__22305),
            .in2(N__17997),
            .in3(N__17833),
            .lcout(\sb_translator_1.state_ledsZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27474),
            .ce(),
            .sr(N__27096));
    defparam \sb_translator_1.send_leds_n_LC_6_8_3 .C_ON=1'b0;
    defparam \sb_translator_1.send_leds_n_LC_6_8_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.send_leds_n_LC_6_8_3 .LUT_INIT=16'b1101110110001100;
    LogicCell40 \sb_translator_1.send_leds_n_LC_6_8_3  (
            .in0(N__17832),
            .in1(N__22062),
            .in2(N__22210),
            .in3(N__27770),
            .lcout(send_leds_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27474),
            .ce(),
            .sr(N__27096));
    defparam \ws2812.new_data_req_RNO_1_LC_6_8_4 .C_ON=1'b0;
    defparam \ws2812.new_data_req_RNO_1_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.new_data_req_RNO_1_LC_6_8_4 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \ws2812.new_data_req_RNO_1_LC_6_8_4  (
            .in0(N__27769),
            .in1(N__25408),
            .in2(_gnd_net_),
            .in3(N__26905),
            .lcout(\ws2812.new_data_req_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_a3_4_LC_6_8_6 .C_ON=1'b0;
    defparam \demux.N_422_i_0_a3_4_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_a3_4_LC_6_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_422_i_0_a3_4_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(N__17380),
            .in2(_gnd_net_),
            .in3(N__23064),
            .lcout(\demux.N_422_i_0_a3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_RNILAHE_10_LC_6_8_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_RNILAHE_10_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_RNILAHE_10_LC_6_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \sb_translator_1.cnt_RNILAHE_10_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(N__17368),
            .in2(_gnd_net_),
            .in3(N__17320),
            .lcout(\sb_translator_1.ram_we_6_0_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_out_2_LC_6_9_0 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_2_LC_6_9_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_2_LC_6_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.instr_out_2_LC_6_9_0  (
            .in0(N__20995),
            .in1(N__21604),
            .in2(N__21575),
            .in3(N__21539),
            .lcout(miso_data_in_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27483),
            .ce(N__23992),
            .sr(N__27102));
    defparam \sb_translator_1.state_RNI2IIJ_0_LC_6_9_1 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNI2IIJ_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNI2IIJ_0_LC_6_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \sb_translator_1.state_RNI2IIJ_0_LC_6_9_1  (
            .in0(N__17235),
            .in1(N__22785),
            .in2(_gnd_net_),
            .in3(N__17050),
            .lcout(\sb_translator_1.num_leds_1_sqmuxa ),
            .ltout(\sb_translator_1.num_leds_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_ram_read_RNO_0_1_LC_6_9_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_ram_read_RNO_0_1_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_ram_read_RNO_0_1_LC_6_9_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \sb_translator_1.cnt_ram_read_RNO_0_1_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__27206),
            .in2(N__17836),
            .in3(N__17831),
            .lcout(\sb_translator_1.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.instr_out_0_LC_6_9_3 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_0_LC_6_9_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_0_LC_6_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.instr_out_0_LC_6_9_3  (
            .in0(N__19971),
            .in1(N__19994),
            .in2(N__19908),
            .in3(N__19930),
            .lcout(miso_data_in_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27483),
            .ce(N__23992),
            .sr(N__27102));
    defparam \sb_translator_1.ram_sel_6_0_0_a2_2_5_LC_6_9_4 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_2_5_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_2_5_LC_6_9_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \sb_translator_1.ram_sel_6_0_0_a2_2_5_LC_6_9_4  (
            .in0(N__17590),
            .in1(N__17642),
            .in2(_gnd_net_),
            .in3(N__17695),
            .lcout(\sb_translator_1.ram_sel_6_0_0_a2_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_sel_6_0_0_a2_3_13_LC_6_9_5 .C_ON=1'b0;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_3_13_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_sel_6_0_0_a2_3_13_LC_6_9_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \sb_translator_1.ram_sel_6_0_0_a2_3_13_LC_6_9_5  (
            .in0(N__17693),
            .in1(N__17643),
            .in2(_gnd_net_),
            .in3(N__17588),
            .lcout(\sb_translator_1.ram_sel_6_0_0_a2_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_0_LC_6_9_6 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_0_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_0_LC_6_9_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \sb_translator_1.ram_we_6_0_0_a2_1_0_LC_6_9_6  (
            .in0(N__17587),
            .in1(N__17641),
            .in2(_gnd_net_),
            .in3(N__17692),
            .lcout(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_3_LC_6_9_7 .C_ON=1'b0;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_3_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.ram_we_6_0_0_a2_1_3_LC_6_9_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \sb_translator_1.ram_we_6_0_0_a2_1_3_LC_6_9_7  (
            .in0(N__17694),
            .in1(N__17644),
            .in2(_gnd_net_),
            .in3(N__17589),
            .lcout(\sb_translator_1.ram_we_6_0_0_a2_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_13_LC_6_10_0 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_13_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_13_LC_6_10_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \demux.N_424_i_0_o2_13_LC_6_10_0  (
            .in0(N__18301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18322),
            .lcout(\demux.N_238 ),
            .ltout(\demux.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_17_LC_6_10_1 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_17_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_17_LC_6_10_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \demux.N_424_i_0_o2_17_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__18273),
            .in2(N__17497),
            .in3(N__18246),
            .lcout(\demux.N_242 ),
            .ltout(\demux.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_34_LC_6_10_2 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_34_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_34_LC_6_10_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \demux.N_424_i_0_a2_34_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__19840),
            .in2(N__17953),
            .in3(N__18356),
            .lcout(\demux.N_424_i_0_a2Z0Z_34 ),
            .ltout(\demux.N_424_i_0_a2Z0Z_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_4_LC_6_10_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_4_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_4_LC_6_10_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \demux.N_424_i_0_a2_4_LC_6_10_3  (
            .in0(N__19810),
            .in1(N__20221),
            .in2(N__17950),
            .in3(N__19756),
            .lcout(\demux.N_424_i_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_LC_6_10_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_LC_6_10_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \demux.N_424_i_0_a2_LC_6_10_4  (
            .in0(N__20319),
            .in1(N__20267),
            .in2(N__20365),
            .in3(N__19666),
            .lcout(\demux.N_424_i_0_aZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_11_LC_6_10_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_11_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_11_LC_6_10_5 .LUT_INIT=16'b1111111011101001;
    LogicCell40 \demux.N_424_i_0_o2_0_11_LC_6_10_5  (
            .in0(N__18357),
            .in1(N__18373),
            .in2(N__20227),
            .in3(N__17905),
            .lcout(\demux.N_424_i_0_o2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_3_LC_6_10_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_3_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_3_LC_6_10_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_424_i_0_o2_0_3_LC_6_10_6  (
            .in0(N__18302),
            .in1(N__18286),
            .in2(N__18253),
            .in3(N__18323),
            .lcout(\demux.N_424_i_0_o2_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_11_LC_6_10_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_11_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_11_LC_6_10_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \demux.N_424_i_0_a2_11_LC_6_10_7  (
            .in0(N__20222),
            .in1(N__19757),
            .in2(N__19818),
            .in3(N__19384),
            .lcout(\demux.N_424_i_0_a2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_1_LC_6_11_0 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_1_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_1_LC_6_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \demux.N_424_i_0_a2_1_LC_6_11_0  (
            .in0(N__18251),
            .in1(N__19532),
            .in2(N__18285),
            .in3(N__18343),
            .lcout(\demux.N_424_i_0_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_38_LC_6_11_1 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_38_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_38_LC_6_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \demux.N_424_i_0_a2_38_LC_6_11_1  (
            .in0(N__17904),
            .in1(N__19844),
            .in2(N__20226),
            .in3(N__18372),
            .lcout(\demux.N_916 ),
            .ltout(\demux.N_916_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_8_LC_6_11_2 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_8_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_8_LC_6_11_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \demux.N_424_i_0_a2_8_LC_6_11_2  (
            .in0(N__19569),
            .in1(N__17880),
            .in2(N__17860),
            .in3(N__17856),
            .lcout(\demux.N_424_i_0_a2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_10_LC_6_11_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_10_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_10_LC_6_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \demux.N_424_i_0_a2_10_LC_6_11_3  (
            .in0(N__18303),
            .in1(N__18341),
            .in2(N__18328),
            .in3(N__19551),
            .lcout(\demux.N_424_i_0_a2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_9_LC_6_11_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_9_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_9_LC_6_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \demux.N_424_i_0_a2_9_LC_6_11_4  (
            .in0(N__18252),
            .in1(N__19533),
            .in2(N__18284),
            .in3(N__18342),
            .lcout(\demux.N_424_i_0_a2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_37_LC_6_11_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_37_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_37_LC_6_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \demux.N_424_i_0_a2_37_LC_6_11_5  (
            .in0(N__20217),
            .in1(N__18371),
            .in2(N__19848),
            .in3(N__18358),
            .lcout(\demux.N_915 ),
            .ltout(\demux.N_915_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_3_LC_6_11_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_3_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_3_LC_6_11_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \demux.N_424_i_0_a2_3_LC_6_11_6  (
            .in0(N__19550),
            .in1(N__18324),
            .in2(N__18307),
            .in3(N__18304),
            .lcout(\demux.N_424_i_0_a2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_12_LC_6_11_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_12_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_12_LC_6_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \demux.N_424_i_0_o2_12_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__18274),
            .in2(_gnd_net_),
            .in3(N__18250),
            .lcout(\demux.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_8_LC_6_12_0 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_8_LC_6_12_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.addr_out_8_LC_6_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_8_LC_6_12_0  (
            .in0(N__21430),
            .in1(N__22198),
            .in2(_gnd_net_),
            .in3(N__19219),
            .lcout(addr_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27500),
            .ce(N__18031),
            .sr(N__27125));
    defparam \sb_translator_1.state_leds_RNIVONR_LC_6_12_1 .C_ON=1'b0;
    defparam \sb_translator_1.state_leds_RNIVONR_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_leds_RNIVONR_LC_6_12_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \sb_translator_1.state_leds_RNIVONR_LC_6_12_1  (
            .in0(N__22197),
            .in1(_gnd_net_),
            .in2(N__17998),
            .in3(N__22873),
            .lcout(\sb_translator_1.state_leds_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_leds_RNIGMAH_LC_6_12_2 .C_ON=1'b0;
    defparam \sb_translator_1.state_leds_RNIGMAH_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_leds_RNIGMAH_LC_6_12_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \sb_translator_1.state_leds_RNIGMAH_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__17993),
            .in2(_gnd_net_),
            .in3(N__22196),
            .lcout(\sb_translator_1.state_leds_RNIGMAHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_13_LC_6_12_3 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_13_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_13_LC_6_12_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \spi_slave_1.miso_RNO_13_LC_6_12_3  (
            .in0(N__17974),
            .in1(N__17968),
            .in2(_gnd_net_),
            .in3(N__18530),
            .lcout(\spi_slave_1.miso_RNOZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_6_LC_6_12_4 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_6_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_6_LC_6_12_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \spi_slave_1.miso_RNO_6_LC_6_12_4  (
            .in0(N__18531),
            .in1(N__18616),
            .in2(_gnd_net_),
            .in3(N__18610),
            .lcout(\spi_slave_1.miso_RNOZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_14_LC_6_12_5 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_14_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_14_LC_6_12_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \spi_slave_1.miso_RNO_14_LC_6_12_5  (
            .in0(N__18595),
            .in1(N__18589),
            .in2(_gnd_net_),
            .in3(N__18581),
            .lcout(),
            .ltout(\spi_slave_1.N_58_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.miso_RNO_9_LC_6_12_6 .C_ON=1'b0;
    defparam \spi_slave_1.miso_RNO_9_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_1.miso_RNO_9_LC_6_12_6 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \spi_slave_1.miso_RNO_9_LC_6_12_6  (
            .in0(N__18532),
            .in1(_gnd_net_),
            .in2(N__18463),
            .in3(N__18460),
            .lcout(\spi_slave_1.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_1.mosi_data_out_15_LC_7_1_5 .C_ON=1'b0;
    defparam \spi_slave_1.mosi_data_out_15_LC_7_1_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_1.mosi_data_out_15_LC_7_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_1.mosi_data_out_15_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18442),
            .lcout(mosi_data_out_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27433),
            .ce(N__18427),
            .sr(N__27069));
    defparam \sb_translator_1.cnt_leds_RNI50UT_5_LC_7_2_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI50UT_5_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI50UT_5_LC_7_2_0 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \sb_translator_1.cnt_leds_RNI50UT_5_LC_7_2_0  (
            .in0(N__18405),
            .in1(N__18858),
            .in2(N__18655),
            .in3(N__20104),
            .lcout(\sb_translator_1.cnt_leds_RNI50UTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIK1VE_5_LC_7_2_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIK1VE_5_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIK1VE_5_LC_7_2_1 .LUT_INIT=16'b1100111100001100;
    LogicCell40 \sb_translator_1.cnt_leds_RNIK1VE_5_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(N__18651),
            .in2(N__18862),
            .in3(N__18403),
            .lcout(\sb_translator_1.cnt_leds_RNIK1VEZ0Z_5 ),
            .ltout(\sb_translator_1.cnt_leds_RNIK1VEZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIB6UT_6_LC_7_2_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIB6UT_6_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIB6UT_6_LC_7_2_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIB6UT_6_LC_7_2_2  (
            .in0(N__18404),
            .in1(N__18832),
            .in2(N__18409),
            .in3(N__18800),
            .lcout(\sb_translator_1.cnt_leds_RNIB6UTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIN4VE_6_LC_7_2_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIN4VE_6_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIN4VE_6_LC_7_2_3 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \sb_translator_1.cnt_leds_RNIN4VE_6_LC_7_2_3  (
            .in0(N__18831),
            .in1(_gnd_net_),
            .in2(N__18804),
            .in3(N__18406),
            .lcout(\sb_translator_1.cnt_leds_RNIN4VEZ0Z_6 ),
            .ltout(\sb_translator_1.cnt_leds_RNIN4VEZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIHCUT_7_LC_7_2_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIHCUT_7_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIHCUT_7_LC_7_2_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIHCUT_7_LC_7_2_4  (
            .in0(N__18765),
            .in1(N__18796),
            .in2(N__18376),
            .in3(N__19245),
            .lcout(\sb_translator_1.cnt_leds_RNIHCUTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIQ7VE_7_LC_7_2_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIQ7VE_7_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIQ7VE_7_LC_7_2_5 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \sb_translator_1.cnt_leds_RNIQ7VE_7_LC_7_2_5  (
            .in0(N__19246),
            .in1(_gnd_net_),
            .in2(N__18805),
            .in3(N__18763),
            .lcout(\sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7 ),
            .ltout(\sb_translator_1.cnt_leds_RNIQ7VEZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNINIUT_8_LC_7_2_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNINIUT_8_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNINIUT_8_LC_7_2_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNINIUT_8_LC_7_2_6  (
            .in0(N__18764),
            .in1(N__18729),
            .in2(N__18769),
            .in3(N__19214),
            .lcout(\sb_translator_1.cnt_leds_RNINIUTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNITAVE_8_LC_7_2_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNITAVE_8_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNITAVE_8_LC_7_2_7 .LUT_INIT=16'b1101010011010100;
    LogicCell40 \sb_translator_1.cnt_leds_RNITAVE_8_LC_7_2_7  (
            .in0(N__19215),
            .in1(N__18766),
            .in2(N__18733),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.cnt_leds_RNITAVEZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_LC_7_3_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIO2NL_0_LC_7_3_0 .LUT_INIT=16'b1110101111010111;
    LogicCell40 \sb_translator_1.cnt_leds_RNIO2NL_0_LC_7_3_0  (
            .in0(N__19097),
            .in1(N__18968),
            .in2(N__19036),
            .in3(N__18995),
            .lcout(\sb_translator_1.N_318_i_i_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIBOUE_2_LC_7_3_1 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIBOUE_2_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIBOUE_2_LC_7_3_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \sb_translator_1.cnt_leds_RNIBOUE_2_LC_7_3_1  (
            .in0(N__18938),
            .in1(N__19073),
            .in2(_gnd_net_),
            .in3(N__19023),
            .lcout(\sb_translator_1.cnt_leds_RNIBOUEZ0Z_2 ),
            .ltout(\sb_translator_1.cnt_leds_RNIBOUEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIPJTT_3_LC_7_3_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIPJTT_3_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIPJTT_3_LC_7_3_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIPJTT_3_LC_7_3_2  (
            .in0(N__19075),
            .in1(N__18910),
            .in2(N__18691),
            .in3(N__18682),
            .lcout(\sb_translator_1.cnt_leds_RNIPJTTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIERUE_3_LC_7_3_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIERUE_3_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIERUE_3_LC_7_3_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \sb_translator_1.cnt_leds_RNIERUE_3_LC_7_3_3  (
            .in0(N__18683),
            .in1(_gnd_net_),
            .in2(N__18916),
            .in3(N__19074),
            .lcout(\sb_translator_1.cnt_leds_RNIERUEZ0Z_3 ),
            .ltout(\sb_translator_1.cnt_leds_RNIERUEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIVPTT_4_LC_7_3_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIVPTT_4_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIVPTT_4_LC_7_3_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIVPTT_4_LC_7_3_4  (
            .in0(N__18650),
            .in1(N__18883),
            .in2(N__18688),
            .in3(N__18681),
            .lcout(\sb_translator_1.cnt_leds_RNIVPTTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIHUUE_4_LC_7_3_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIHUUE_4_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIHUUE_4_LC_7_3_5 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \sb_translator_1.cnt_leds_RNIHUUE_4_LC_7_3_5  (
            .in0(N__18684),
            .in1(_gnd_net_),
            .in2(N__18889),
            .in3(N__18649),
            .lcout(\sb_translator_1.cnt_leds_RNIHUUEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI8LUE_1_LC_7_3_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI8LUE_1_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI8LUE_1_LC_7_3_6 .LUT_INIT=16'b1011001010110010;
    LogicCell40 \sb_translator_1.cnt_leds_RNI8LUE_1_LC_7_3_6  (
            .in0(N__19096),
            .in1(N__18967),
            .in2(N__19035),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.state56_a_5_44 ),
            .ltout(\sb_translator_1.state56_a_5_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIJDTT_2_LC_7_3_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIJDTT_2_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIJDTT_2_LC_7_3_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIJDTT_2_LC_7_3_7  (
            .in0(N__18937),
            .in1(N__19072),
            .in2(N__19045),
            .in3(N__19019),
            .lcout(\sb_translator_1.cnt_leds_RNIJDTTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_0_LC_7_4_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_0_LC_7_4_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_0_LC_7_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_0_LC_7_4_0  (
            .in0(N__22323),
            .in1(N__18996),
            .in2(_gnd_net_),
            .in3(N__18973),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(\sb_translator_1.cnt_leds_cry_0 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_1_LC_7_4_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_1_LC_7_4_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_1_LC_7_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_1_LC_7_4_1  (
            .in0(N__22334),
            .in1(N__18969),
            .in2(_gnd_net_),
            .in3(N__18943),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_1 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_0 ),
            .carryout(\sb_translator_1.cnt_leds_cry_1 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_2_LC_7_4_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_2_LC_7_4_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_2_LC_7_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_2_LC_7_4_2  (
            .in0(N__22324),
            .in1(N__18939),
            .in2(_gnd_net_),
            .in3(N__18919),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_2 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_1 ),
            .carryout(\sb_translator_1.cnt_leds_cry_2 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_3_LC_7_4_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_3_LC_7_4_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_3_LC_7_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_3_LC_7_4_3  (
            .in0(N__22335),
            .in1(N__18914),
            .in2(_gnd_net_),
            .in3(N__18892),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_3 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_2 ),
            .carryout(\sb_translator_1.cnt_leds_cry_3 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_4_LC_7_4_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_4_LC_7_4_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_4_LC_7_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_4_LC_7_4_4  (
            .in0(N__22325),
            .in1(N__18887),
            .in2(_gnd_net_),
            .in3(N__18865),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_4 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_3 ),
            .carryout(\sb_translator_1.cnt_leds_cry_4 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_5_LC_7_4_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_5_LC_7_4_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_5_LC_7_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_5_LC_7_4_5  (
            .in0(N__22336),
            .in1(N__18856),
            .in2(_gnd_net_),
            .in3(N__18835),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_5 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_4 ),
            .carryout(\sb_translator_1.cnt_leds_cry_5 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_6_LC_7_4_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_6_LC_7_4_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_6_LC_7_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_6_LC_7_4_6  (
            .in0(N__22326),
            .in1(N__18829),
            .in2(_gnd_net_),
            .in3(N__18808),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_6 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_5 ),
            .carryout(\sb_translator_1.cnt_leds_cry_6 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_7_LC_7_4_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_7_LC_7_4_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_7_LC_7_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_7_LC_7_4_7  (
            .in0(N__22337),
            .in1(N__19243),
            .in2(_gnd_net_),
            .in3(N__19222),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_7 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_6 ),
            .carryout(\sb_translator_1.cnt_leds_cry_7 ),
            .clk(N__27453),
            .ce(N__19355),
            .sr(N__27081));
    defparam \sb_translator_1.cnt_leds_8_LC_7_5_0 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_8_LC_7_5_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_8_LC_7_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_8_LC_7_5_0  (
            .in0(N__22333),
            .in1(N__19213),
            .in2(_gnd_net_),
            .in3(N__19192),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\sb_translator_1.cnt_leds_cry_8 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_9_LC_7_5_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_9_LC_7_5_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_9_LC_7_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_9_LC_7_5_1  (
            .in0(N__22321),
            .in1(N__21352),
            .in2(_gnd_net_),
            .in3(N__19189),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_9 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_8 ),
            .carryout(\sb_translator_1.cnt_leds_cry_9 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_10_LC_7_5_2 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_10_LC_7_5_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_10_LC_7_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_10_LC_7_5_2  (
            .in0(N__22330),
            .in1(N__19186),
            .in2(_gnd_net_),
            .in3(N__19156),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_10 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_9 ),
            .carryout(\sb_translator_1.cnt_leds_cry_10 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_11_LC_7_5_3 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_11_LC_7_5_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_11_LC_7_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_11_LC_7_5_3  (
            .in0(N__22318),
            .in1(N__19151),
            .in2(_gnd_net_),
            .in3(N__19120),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_11 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_10 ),
            .carryout(\sb_translator_1.cnt_leds_cry_11 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_12_LC_7_5_4 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_12_LC_7_5_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_12_LC_7_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_12_LC_7_5_4  (
            .in0(N__22331),
            .in1(N__21391),
            .in2(_gnd_net_),
            .in3(N__19117),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_12 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_11 ),
            .carryout(\sb_translator_1.cnt_leds_cry_12 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_13_LC_7_5_5 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_13_LC_7_5_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_13_LC_7_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_13_LC_7_5_5  (
            .in0(N__22319),
            .in1(N__20842),
            .in2(_gnd_net_),
            .in3(N__19114),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_13 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_12 ),
            .carryout(\sb_translator_1.cnt_leds_cry_13 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_14_LC_7_5_6 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_14_LC_7_5_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_14_LC_7_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_14_LC_7_5_6  (
            .in0(N__22332),
            .in1(N__20743),
            .in2(_gnd_net_),
            .in3(N__19111),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_14 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_13 ),
            .carryout(\sb_translator_1.cnt_leds_cry_14 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_15_LC_7_5_7 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_15_LC_7_5_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_15_LC_7_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \sb_translator_1.cnt_leds_15_LC_7_5_7  (
            .in0(N__22320),
            .in1(N__20905),
            .in2(_gnd_net_),
            .in3(N__19372),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_15 ),
            .ltout(),
            .carryin(\sb_translator_1.cnt_leds_cry_14 ),
            .carryout(\sb_translator_1.cnt_leds_cry_15 ),
            .clk(N__27460),
            .ce(N__19366),
            .sr(N__27086));
    defparam \sb_translator_1.cnt_leds_16_LC_7_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_16_LC_7_6_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.cnt_leds_16_LC_7_6_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \sb_translator_1.cnt_leds_16_LC_7_6_0  (
            .in0(N__20599),
            .in1(N__22322),
            .in2(_gnd_net_),
            .in3(N__19369),
            .lcout(\sb_translator_1.cnt_ledsZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27468),
            .ce(N__19365),
            .sr(N__27091));
    defparam \sb_translator_1.rgb_data_tmp_2_LC_7_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_2_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_2_LC_7_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_2_LC_7_7_0  (
            .in0(N__20980),
            .in1(N__21619),
            .in2(N__21574),
            .in3(N__21538),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27475),
            .ce(N__25430),
            .sr(N__27097));
    defparam \demux.N_424_i_0_a3_4_LC_7_7_2 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a3_4_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a3_4_LC_7_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_424_i_0_a3_4_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__23073),
            .lcout(\demux.N_424_i_0_a3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_1_LC_7_7_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_1_LC_7_7_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \demux.N_424_i_0_o2_1_LC_7_7_3  (
            .in0(N__19327),
            .in1(N__23371),
            .in2(_gnd_net_),
            .in3(N__20644),
            .lcout(),
            .ltout(\demux.N_424_i_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_7_LC_7_7_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_7_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_7_LC_7_7_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \demux.N_424_i_0_o2_7_LC_7_7_4  (
            .in0(N__19315),
            .in1(N__19309),
            .in2(N__19294),
            .in3(N__23302),
            .lcout(\demux.N_424_i_0_o2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a3_LC_7_7_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a3_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a3_LC_7_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_424_i_0_a3_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__19291),
            .in2(_gnd_net_),
            .in3(N__25836),
            .lcout(\demux.N_424_i_0_aZ0Z3 ),
            .ltout(\demux.N_424_i_0_aZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_0_LC_7_7_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_0_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_0_LC_7_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_0_LC_7_7_6  (
            .in0(N__20001),
            .in1(N__19947),
            .in2(N__19276),
            .in3(N__19894),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27475),
            .ce(N__25430),
            .sr(N__27097));
    defparam \demux.N_421_i_0_o2_0_LC_7_8_1 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_0_LC_7_8_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_421_i_0_o2_0_LC_7_8_1  (
            .in0(N__23477),
            .in1(N__19273),
            .in2(N__19261),
            .in3(N__23408),
            .lcout(),
            .ltout(\demux.N_421_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_2_LC_7_8_2 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_2_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_2_LC_7_8_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_421_i_0_o2_2_LC_7_8_2  (
            .in0(N__19519),
            .in1(N__23367),
            .in2(N__19507),
            .in3(N__19390),
            .lcout(\demux.N_421_i_0_o2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_a3_LC_7_8_3 .C_ON=1'b0;
    defparam \demux.N_422_i_0_a3_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_a3_LC_7_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \demux.N_422_i_0_a3_LC_7_8_3  (
            .in0(N__25837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19504),
            .lcout(\demux.N_422_i_0_aZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_0_LC_7_8_4 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_0_LC_7_8_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \demux.N_422_i_0_o2_0_LC_7_8_4  (
            .in0(N__19489),
            .in1(N__19477),
            .in2(N__23424),
            .in3(N__23478),
            .lcout(),
            .ltout(\demux.N_422_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_1_LC_7_8_5 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_1_LC_7_8_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \demux.N_422_i_0_o2_1_LC_7_8_5  (
            .in0(N__23368),
            .in1(_gnd_net_),
            .in2(N__19465),
            .in3(N__19462),
            .lcout(),
            .ltout(\demux.N_422_i_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_7_LC_7_8_6 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_7_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_7_LC_7_8_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \demux.N_422_i_0_o2_7_LC_7_8_6  (
            .in0(N__19450),
            .in1(N__19444),
            .in2(N__19432),
            .in3(N__23298),
            .lcout(\demux.N_422_i_0_o2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_a3_5_LC_7_9_0 .C_ON=1'b0;
    defparam \demux.N_423_i_0_a3_5_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_a3_5_LC_7_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_423_i_0_a3_5_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__23297),
            .in2(_gnd_net_),
            .in3(N__19429),
            .lcout(),
            .ltout(\demux.N_423_i_0_a3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_2_LC_7_9_1 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_2_LC_7_9_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_423_i_0_o2_2_LC_7_9_1  (
            .in0(N__19417),
            .in1(N__23346),
            .in2(N__19405),
            .in3(N__19672),
            .lcout(\demux.N_423_i_0_o2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_a3_4_LC_7_9_2 .C_ON=1'b0;
    defparam \demux.N_421_i_0_a3_4_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_a3_4_LC_7_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_421_i_0_a3_4_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__23055),
            .in2(_gnd_net_),
            .in3(N__19402),
            .lcout(\demux.N_837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_12_LC_7_9_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_12_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_12_LC_7_9_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \demux.N_424_i_0_a2_12_LC_7_9_3  (
            .in0(N__19817),
            .in1(N__19767),
            .in2(_gnd_net_),
            .in3(N__19383),
            .lcout(\demux.N_918 ),
            .ltout(\demux.N_918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_5_LC_7_9_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_5_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_5_LC_7_9_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \demux.N_424_i_0_a2_5_LC_7_9_4  (
            .in0(N__20316),
            .in1(N__20361),
            .in2(N__19705),
            .in3(N__20274),
            .lcout(\demux.N_424_i_0_a2Z0Z_5 ),
            .ltout(\demux.N_424_i_0_a2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_0_LC_7_9_5 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_0_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_0_LC_7_9_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_423_i_0_o2_0_LC_7_9_5  (
            .in0(N__23452),
            .in1(N__19702),
            .in2(N__19690),
            .in3(N__19687),
            .lcout(\demux.N_423_i_0_o2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_7_LC_7_9_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_7_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_7_LC_7_9_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \demux.N_424_i_0_a2_7_LC_7_9_6  (
            .in0(N__20318),
            .in1(N__20359),
            .in2(N__20275),
            .in3(N__19665),
            .lcout(\demux.N_424_i_0_a2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_44_LC_7_9_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_44_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_44_LC_7_9_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \demux.N_424_i_0_a2_44_LC_7_9_7  (
            .in0(N__20360),
            .in1(N__20273),
            .in2(_gnd_net_),
            .in3(N__20317),
            .lcout(\demux.N_917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_13_LC_7_10_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_13_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_13_LC_7_10_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_13_LC_7_10_1  (
            .in0(N__25848),
            .in1(N__25747),
            .in2(N__25723),
            .in3(N__25655),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27496),
            .ce(N__21503),
            .sr(N__27115));
    defparam \sb_translator_1.rgb_data_tmp_11_LC_7_10_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_11_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_11_LC_7_10_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \sb_translator_1.rgb_data_tmp_11_LC_7_10_2  (
            .in0(N__24220),
            .in1(N__25849),
            .in2(N__24263),
            .in3(N__24177),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27496),
            .ce(N__21503),
            .sr(N__27115));
    defparam \demux.N_424_i_0_o2_0_8_1_LC_7_10_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_8_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_8_1_LC_7_10_3 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \demux.N_424_i_0_o2_0_8_1_LC_7_10_3  (
            .in0(N__19615),
            .in1(N__19603),
            .in2(_gnd_net_),
            .in3(N__19576),
            .lcout(),
            .ltout(\demux.N_424_i_0_o2_0_8Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_8_LC_7_10_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_8_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_8_LC_7_10_4 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \demux.N_424_i_0_o2_0_8_LC_7_10_4  (
            .in0(N__19558),
            .in1(N__19552),
            .in2(N__19537),
            .in3(N__19534),
            .lcout(),
            .ltout(\demux.N_424_i_0_o2_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_LC_7_10_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_LC_7_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \demux.N_424_i_0_o2_0_LC_7_10_5  (
            .in0(N__19729),
            .in1(N__20062),
            .in2(N__20056),
            .in3(N__20053),
            .lcout(\demux.N_424_i_0_o2Z0Z_0 ),
            .ltout(\demux.N_424_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_9_LC_7_10_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_9_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_9_LC_7_10_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_9_LC_7_10_6  (
            .in0(N__24092),
            .in1(N__24121),
            .in2(N__20047),
            .in3(N__24044),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27496),
            .ce(N__21503),
            .sr(N__27115));
    defparam \demux.N_424_i_0_o2_4_LC_7_11_0 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_4_LC_7_11_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_424_i_0_o2_4_LC_7_11_0  (
            .in0(N__20044),
            .in1(N__24478),
            .in2(N__20032),
            .in3(N__24411),
            .lcout(),
            .ltout(\demux.N_424_i_0_o2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_8_LC_7_11_1 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_8_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_8_LC_7_11_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_424_i_0_o2_8_LC_7_11_1  (
            .in0(N__24326),
            .in1(N__20017),
            .in2(N__20005),
            .in3(N__19858),
            .lcout(\demux.N_424_i_0_o2Z0Z_8 ),
            .ltout(\demux.N_424_i_0_o2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_8_LC_7_11_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_8_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_8_LC_7_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_8_LC_7_11_2  (
            .in0(N__19975),
            .in1(N__19948),
            .in2(N__19912),
            .in3(N__19909),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27501),
            .ce(N__21517),
            .sr(N__27126));
    defparam \demux.N_424_i_0_a3_7_LC_7_11_3 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a3_7_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a3_7_LC_7_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \demux.N_424_i_0_a3_7_LC_7_11_3  (
            .in0(N__23931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19876),
            .lcout(\demux.N_424_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_a2_33_LC_7_11_4 .C_ON=1'b0;
    defparam \demux.N_424_i_0_a2_33_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_a2_33_LC_7_11_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \demux.N_424_i_0_a2_33_LC_7_11_4  (
            .in0(N__20269),
            .in1(_gnd_net_),
            .in2(N__20320),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\demux.N_906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_4_LC_7_11_5 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_4_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_4_LC_7_11_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \demux.N_424_i_0_o2_0_4_LC_7_11_5  (
            .in0(N__19852),
            .in1(N__19819),
            .in2(N__19771),
            .in3(N__19768),
            .lcout(\demux.N_424_i_0_o2_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_a3_7_LC_7_11_6 .C_ON=1'b0;
    defparam \demux.N_420_i_0_a3_7_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_a3_7_LC_7_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_420_i_0_a3_7_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__19723),
            .in2(_gnd_net_),
            .in3(N__23930),
            .lcout(\demux.N_420_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_15_LC_7_11_7 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_15_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_15_LC_7_11_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \demux.N_424_i_0_o2_15_LC_7_11_7  (
            .in0(N__20358),
            .in1(N__20312),
            .in2(_gnd_net_),
            .in3(N__20268),
            .lcout(\demux.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_a3_7_LC_7_12_7 .C_ON=1'b0;
    defparam \demux.N_419_i_0_a3_7_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_a3_7_LC_7_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_419_i_0_a3_7_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__23922),
            .in2(_gnd_net_),
            .in3(N__20197),
            .lcout(\demux.N_419_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_0_c_THRU_CRY_0_LC_8_3_0 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_0_c_THRU_CRY_0_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_0_c_THRU_CRY_0_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \sb_translator_1.state56_a_5_cry_0_c_THRU_CRY_0_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__20172),
            .in2(N__20179),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\sb_translator_1.state56_a_5_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIJ5J22_0_LC_8_3_1 .C_ON=1'b1;
    defparam \sb_translator_1.cnt_leds_RNIJ5J22_0_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIJ5J22_0_LC_8_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.cnt_leds_RNIJ5J22_0_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__20158),
            .in2(N__20152),
            .in3(N__20143),
            .lcout(\sb_translator_1.state56_a_5_2 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_0_c_THRU_CO ),
            .carryout(\sb_translator_1.state56_a_5_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_0_c_RNIUH4N1_LC_8_3_2 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_0_c_RNIUH4N1_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_0_c_RNIUH4N1_LC_8_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_0_c_RNIUH4N1_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__20140),
            .in2(N__20134),
            .in3(N__20125),
            .lcout(\sb_translator_1.state56_a_5_3 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_0 ),
            .carryout(\sb_translator_1.state56_a_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_1_c_RNI8T5N1_LC_8_3_3 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_1_c_RNI8T5N1_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_1_c_RNI8T5N1_LC_8_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_1_c_RNI8T5N1_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__20122),
            .in2(N__20116),
            .in3(N__20107),
            .lcout(\sb_translator_1.state56_a_5_4 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_1 ),
            .carryout(\sb_translator_1.state56_a_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNII87N1_LC_8_3_4 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNII87N1_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNII87N1_LC_8_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_2_c_RNII87N1_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__20103),
            .in2(N__20092),
            .in3(N__20083),
            .lcout(\sb_translator_1.state56_a_5_5 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_2 ),
            .carryout(\sb_translator_1.state56_a_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_3_c_RNISJ8N1_LC_8_3_5 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_3_c_RNISJ8N1_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_3_c_RNISJ8N1_LC_8_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_3_c_RNISJ8N1_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__20080),
            .in2(N__20074),
            .in3(N__20065),
            .lcout(\sb_translator_1.state56_a_5_6 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_3 ),
            .carryout(\sb_translator_1.state56_a_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_4_c_RNI6V9N1_LC_8_3_6 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_4_c_RNI6V9N1_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_4_c_RNI6V9N1_LC_8_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_4_c_RNI6V9N1_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__20521),
            .in2(N__20515),
            .in3(N__20506),
            .lcout(\sb_translator_1.state56_a_5_7 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_4 ),
            .carryout(\sb_translator_1.state56_a_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_5_c_RNIGABN1_LC_8_3_7 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_5_c_RNIGABN1_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_5_c_RNIGABN1_LC_8_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_5_c_RNIGABN1_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__20503),
            .in2(N__20497),
            .in3(N__20488),
            .lcout(\sb_translator_1.state56_a_5_8 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_5 ),
            .carryout(\sb_translator_1.state56_a_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_6_c_RNIQLCN1_LC_8_4_0 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_6_c_RNIQLCN1_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_6_c_RNIQLCN1_LC_8_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_6_c_RNIQLCN1_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__20485),
            .in2(N__20475),
            .in3(N__20452),
            .lcout(\sb_translator_1.state56_a_5_9 ),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\sb_translator_1.state56_a_5_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_7_c_RNII4T22_LC_8_4_1 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_7_c_RNII4T22_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_7_c_RNII4T22_LC_8_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_7_c_RNII4T22_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(N__20440),
            .in3(N__20422),
            .lcout(\sb_translator_1.state56_a_5_10 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_7 ),
            .carryout(\sb_translator_1.state56_a_5_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_8_c_RNIVTUS2_LC_8_4_2 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_8_c_RNIVTUS2_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_8_c_RNIVTUS2_LC_8_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_8_c_RNIVTUS2_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__20419),
            .in2(N__20410),
            .in3(N__20398),
            .lcout(\sb_translator_1.state56_a_5_11 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_8 ),
            .carryout(\sb_translator_1.state56_a_5_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_9_c_RNINN433_LC_8_4_3 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_9_c_RNINN433_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_9_c_RNINN433_LC_8_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_9_c_RNINN433_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__20395),
            .in2(N__20386),
            .in3(N__20374),
            .lcout(\sb_translator_1.state56_a_5_12 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_9 ),
            .carryout(\sb_translator_1.state56_a_5_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNI8BIQ2_LC_8_4_4 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNI8BIQ2_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNI8BIQ2_LC_8_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_10_c_RNI8BIQ2_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__20554),
            .in2(N__20574),
            .in3(N__20371),
            .lcout(\sb_translator_1.state56_a_5_13 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_10 ),
            .carryout(\sb_translator_1.state56_a_5_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_11_c_RNIIMJQ2_LC_8_4_5 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_11_c_RNIIMJQ2_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_11_c_RNIIMJQ2_LC_8_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_11_c_RNIIMJQ2_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__20827),
            .in2(N__20728),
            .in3(N__20368),
            .lcout(\sb_translator_1.state56_a_5_14 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_11 ),
            .carryout(\sb_translator_1.state56_a_5_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIS1LQ2_LC_8_4_6 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIS1LQ2_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIS1LQ2_LC_8_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_12_c_RNIS1LQ2_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(N__20530),
            .in2(N__20545),
            .in3(N__20608),
            .lcout(\sb_translator_1.state56_a_5_15 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_12 ),
            .carryout(\sb_translator_1.state56_a_5_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNIK1552_LC_8_4_7 .C_ON=1'b1;
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNIK1552_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNIK1552_LC_8_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \sb_translator_1.state56_a_5_cry_13_c_RNIK1552_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(N__20584),
            .in2(N__20890),
            .in3(N__20605),
            .lcout(\sb_translator_1.state56_a_5_16 ),
            .ltout(),
            .carryin(\sb_translator_1.state56_a_5_cry_13 ),
            .carryout(\sb_translator_1.state56_a_5_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_14_c_RNI7UEO_LC_8_5_0 .C_ON=1'b0;
    defparam \sb_translator_1.state56_a_5_cry_14_c_RNI7UEO_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_14_c_RNI7UEO_LC_8_5_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \sb_translator_1.state56_a_5_cry_14_c_RNI7UEO_LC_8_5_0  (
            .in0(N__20916),
            .in1(N__20949),
            .in2(_gnd_net_),
            .in3(N__20602),
            .lcout(\sb_translator_1.state56_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_15_LC_8_5_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_15_LC_8_5_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.num_leds_15_LC_8_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.num_leds_15_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22945),
            .lcout(\sb_translator_1.num_ledsZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27469),
            .ce(N__22355),
            .sr(N__27092));
    defparam \sb_translator_1.cnt_leds_RNI7Q5F_16_LC_8_6_0 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI7Q5F_16_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI7Q5F_16_LC_8_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \sb_translator_1.cnt_leds_RNI7Q5F_16_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20598),
            .lcout(\sb_translator_1.cnt_leds_i_16 ),
            .ltout(\sb_translator_1.cnt_leds_i_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.num_leds_RNIOJBM_15_LC_8_6_1 .C_ON=1'b0;
    defparam \sb_translator_1.num_leds_RNIOJBM_15_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.num_leds_RNIOJBM_15_LC_8_6_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \sb_translator_1.num_leds_RNIOJBM_15_LC_8_6_1  (
            .in0(N__20947),
            .in1(_gnd_net_),
            .in2(N__20587),
            .in3(_gnd_net_),
            .lcout(\sb_translator_1.num_leds_RNIOJBMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIV62R1_13_LC_8_6_2 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIV62R1_13_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIV62R1_13_LC_8_6_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \sb_translator_1.cnt_leds_RNIV62R1_13_LC_8_6_2  (
            .in0(N__20575),
            .in1(N__20877),
            .in2(N__20782),
            .in3(N__20840),
            .lcout(\sb_translator_1.cnt_leds_RNIV62R1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI48HT_14_LC_8_6_3 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI48HT_14_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI48HT_14_LC_8_6_3 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \sb_translator_1.cnt_leds_RNI48HT_14_LC_8_6_3  (
            .in0(N__20812),
            .in1(N__20781),
            .in2(_gnd_net_),
            .in3(N__20742),
            .lcout(\sb_translator_1.cnt_leds_RNI48HTZ0Z_14 ),
            .ltout(\sb_translator_1.cnt_leds_RNI48HTZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIBJ2R1_15_LC_8_6_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIBJ2R1_15_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIBJ2R1_15_LC_8_6_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNIBJ2R1_15_LC_8_6_4  (
            .in0(N__20903),
            .in1(N__20946),
            .in2(N__20533),
            .in3(N__20814),
            .lcout(\sb_translator_1.cnt_leds_RNIBJ2R1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNIE5NC1_15_LC_8_6_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNIE5NC1_15_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNIE5NC1_15_LC_8_6_5 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \sb_translator_1.cnt_leds_RNIE5NC1_15_LC_8_6_5  (
            .in0(N__20815),
            .in1(N__20948),
            .in2(N__20920),
            .in3(N__20904),
            .lcout(\sb_translator_1.cnt_leds_RNIE5NC1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI15HT_13_LC_8_6_6 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI15HT_13_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI15HT_13_LC_8_6_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \sb_translator_1.cnt_leds_RNI15HT_13_LC_8_6_6  (
            .in0(N__20780),
            .in1(N__20878),
            .in2(_gnd_net_),
            .in3(N__20841),
            .lcout(\sb_translator_1.cnt_leds_RNI15HTZ0Z_13 ),
            .ltout(\sb_translator_1.cnt_leds_RNI15HTZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI5D2R1_14_LC_8_6_7 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI5D2R1_14_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI5D2R1_14_LC_8_6_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \sb_translator_1.cnt_leds_RNI5D2R1_14_LC_8_6_7  (
            .in0(N__20813),
            .in1(N__20776),
            .in2(N__20746),
            .in3(N__20741),
            .lcout(\sb_translator_1.cnt_leds_RNI5D2R1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_8_LC_8_7_1 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_8_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_8_LC_8_7_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \demux.N_422_i_0_o2_8_LC_8_7_1  (
            .in0(N__23809),
            .in1(N__24361),
            .in2(N__20716),
            .in3(N__21268),
            .lcout(\demux.N_422_i_0_o2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_4_LC_8_7_4 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_4_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_4_LC_8_7_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_418_i_0_o2_4_LC_8_7_4  (
            .in0(N__20701),
            .in1(N__24435),
            .in2(N__20686),
            .in3(N__23956),
            .lcout(\demux.N_418_i_0_o2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_424_i_0_o2_0_0_LC_8_7_6 .C_ON=1'b0;
    defparam \demux.N_424_i_0_o2_0_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_424_i_0_o2_0_0_LC_8_7_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_424_i_0_o2_0_0_LC_8_7_6  (
            .in0(N__23479),
            .in1(N__20674),
            .in2(N__20659),
            .in3(N__23412),
            .lcout(\demux.N_424_i_0_o2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_a3_4_LC_8_7_7 .C_ON=1'b0;
    defparam \demux.N_420_i_0_a3_4_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_a3_4_LC_8_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_420_i_0_a3_4_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__20638),
            .in2(_gnd_net_),
            .in3(N__23074),
            .lcout(\demux.N_420_i_0_a3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_a3_9_LC_8_8_0 .C_ON=1'b0;
    defparam \demux.N_418_i_0_a3_9_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_a3_9_LC_8_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_418_i_0_a3_9_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__20623),
            .in2(_gnd_net_),
            .in3(N__24505),
            .lcout(),
            .ltout(\demux.N_884_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_8_LC_8_8_1 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_8_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_8_LC_8_8_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \demux.N_418_i_0_o2_8_LC_8_8_1  (
            .in0(N__21154),
            .in1(N__21148),
            .in2(N__21133),
            .in3(N__21073),
            .lcout(\demux.N_418_i_0_o2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_a3_7_LC_8_8_3 .C_ON=1'b0;
    defparam \demux.N_421_i_0_a3_7_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_a3_7_LC_8_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_421_i_0_a3_7_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__23951),
            .in2(_gnd_net_),
            .in3(N__21130),
            .lcout(\demux.N_421_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_4_LC_8_8_4 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_4_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_4_LC_8_8_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_421_i_0_o2_4_LC_8_8_4  (
            .in0(N__21115),
            .in1(N__24504),
            .in2(N__21100),
            .in3(N__24434),
            .lcout(),
            .ltout(\demux.N_421_i_0_o2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_8_LC_8_8_5 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_8_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_8_LC_8_8_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_421_i_0_o2_8_LC_8_8_5  (
            .in0(N__21088),
            .in1(N__21072),
            .in2(N__21025),
            .in3(N__21022),
            .lcout(),
            .ltout(\demux.N_421_i_0_o2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_421_i_0_o2_10_LC_8_8_6 .C_ON=1'b0;
    defparam \demux.N_421_i_0_o2_10_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_421_i_0_o2_10_LC_8_8_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_421_i_0_o2_10_LC_8_8_6  (
            .in0(N__21016),
            .in1(N__23296),
            .in2(N__21004),
            .in3(N__21001),
            .lcout(\demux.N_421_i_0_o2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_15_LC_8_9_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_15_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_15_LC_8_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_15_LC_8_9_0  (
            .in0(N__23714),
            .in1(N__23884),
            .in2(N__23700),
            .in3(N__23771),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27497),
            .ce(N__21516),
            .sr(N__27116));
    defparam \sb_translator_1.rgb_data_tmp_14_LC_8_9_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_14_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_14_LC_8_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_14_LC_8_9_1  (
            .in0(N__23617),
            .in1(N__23645),
            .in2(N__23588),
            .in3(N__23558),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27497),
            .ce(N__21516),
            .sr(N__27116));
    defparam \sb_translator_1.rgb_data_tmp_12_LC_8_9_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_12_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_12_LC_8_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_12_LC_8_9_2  (
            .in0(N__25623),
            .in1(N__25574),
            .in2(N__25539),
            .in3(N__25477),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27497),
            .ce(N__21516),
            .sr(N__27116));
    defparam \sb_translator_1.rgb_data_tmp_10_LC_8_9_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_10_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_10_LC_8_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_10_LC_8_9_3  (
            .in0(N__20990),
            .in1(N__21614),
            .in2(N__21583),
            .in3(N__21540),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27497),
            .ce(N__21516),
            .sr(N__27116));
    defparam \sb_translator_1.addr_out_RNO_0_8_LC_8_9_4 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_8_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_8_LC_8_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_8_LC_8_9_4  (
            .in0(N__23008),
            .in1(N__21469),
            .in2(_gnd_net_),
            .in3(N__21457),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_2_9_LC_8_9_5 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_2_9_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI1VFQ_2_9_LC_8_9_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \sb_translator_1.cnt_leds_RNI1VFQ_2_9_LC_8_9_5  (
            .in0(N__21997),
            .in1(N__21416),
            .in2(_gnd_net_),
            .in3(N__21363),
            .lcout(\sb_translator_1.cnt_leds_RNI1VFQ_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_a3_7_LC_8_10_0 .C_ON=1'b0;
    defparam \demux.N_422_i_0_a3_7_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_a3_7_LC_8_10_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \demux.N_422_i_0_a3_7_LC_8_10_0  (
            .in0(N__23950),
            .in1(_gnd_net_),
            .in2(N__21283),
            .in3(_gnd_net_),
            .lcout(\demux.N_422_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_7_LC_8_10_1 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_7_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_7_LC_8_10_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_417_i_0_o2_7_LC_8_10_1  (
            .in0(N__23295),
            .in1(N__21259),
            .in2(N__21739),
            .in3(N__21760),
            .lcout(\demux.N_417_i_0_o2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_a3_7_LC_8_10_3 .C_ON=1'b0;
    defparam \demux.N_423_i_0_a3_7_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_a3_7_LC_8_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_423_i_0_a3_7_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__23949),
            .in2(_gnd_net_),
            .in3(N__21247),
            .lcout(\demux.N_423_i_0_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_4_LC_8_10_4 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_4_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_4_LC_8_10_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_423_i_0_o2_4_LC_8_10_4  (
            .in0(N__21229),
            .in1(N__24506),
            .in2(N__21217),
            .in3(N__24436),
            .lcout(),
            .ltout(\demux.N_423_i_0_o2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_8_LC_8_10_5 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_8_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_8_LC_8_10_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_423_i_0_o2_8_LC_8_10_5  (
            .in0(N__21202),
            .in1(N__24354),
            .in2(N__21187),
            .in3(N__21184),
            .lcout(),
            .ltout(\demux.N_423_i_0_o2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_423_i_0_o2_10_LC_8_10_6 .C_ON=1'b0;
    defparam \demux.N_423_i_0_o2_10_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_423_i_0_o2_10_LC_8_10_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_423_i_0_o2_10_LC_8_10_6  (
            .in0(N__21178),
            .in1(N__23072),
            .in2(N__21163),
            .in3(N__21160),
            .lcout(\demux.N_423_i_0_o2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_0_LC_8_11_0 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_0_LC_8_11_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_417_i_0_o2_0_LC_8_11_0  (
            .in0(N__23480),
            .in1(N__21808),
            .in2(N__23425),
            .in3(N__21796),
            .lcout(),
            .ltout(\demux.N_417_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_1_LC_8_11_1 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_1_LC_8_11_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \demux.N_417_i_0_o2_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__21778),
            .in2(N__21763),
            .in3(N__23369),
            .lcout(\demux.N_417_i_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_a3_4_LC_8_11_3 .C_ON=1'b0;
    defparam \demux.N_417_i_0_a3_4_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_a3_4_LC_8_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_417_i_0_a3_4_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__21754),
            .in2(_gnd_net_),
            .in3(N__23056),
            .lcout(\demux.N_417_i_0_a3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_0_LC_8_11_4 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_0_LC_8_11_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_419_i_0_o2_0_LC_8_11_4  (
            .in0(N__23481),
            .in1(N__21730),
            .in2(N__23426),
            .in3(N__21718),
            .lcout(),
            .ltout(\demux.N_419_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_2_LC_8_11_5 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_2_LC_8_11_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_419_i_0_o2_2_LC_8_11_5  (
            .in0(N__21700),
            .in1(N__23370),
            .in2(N__21685),
            .in3(N__21655),
            .lcout(),
            .ltout(\demux.N_419_i_0_o2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_10_LC_8_11_6 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_10_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_10_LC_8_11_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_419_i_0_o2_10_LC_8_11_6  (
            .in0(N__23057),
            .in1(N__21682),
            .in2(N__21667),
            .in3(N__21625),
            .lcout(\demux.N_419_i_0_o2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_a3_5_LC_8_11_7 .C_ON=1'b0;
    defparam \demux.N_419_i_0_a3_5_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_a3_5_LC_8_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_419_i_0_a3_5_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__23272),
            .in2(_gnd_net_),
            .in3(N__21664),
            .lcout(\demux.N_419_i_0_a3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_8_LC_8_12_6 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_8_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_8_LC_8_12_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \demux.N_419_i_0_o2_8_LC_8_12_6  (
            .in0(N__24353),
            .in1(N__24526),
            .in2(N__21649),
            .in3(N__21631),
            .lcout(\demux.N_419_i_0_o2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNILP7UD_LC_9_3_0 .C_ON=1'b0;
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNILP7UD_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_2_c_RNILP7UD_LC_9_3_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \sb_translator_1.state56_a_5_cry_2_c_RNILP7UD_LC_9_3_0  (
            .in0(N__22471),
            .in1(N__22465),
            .in2(N__22459),
            .in3(N__22105),
            .lcout(),
            .ltout(\sb_translator_1.N_318_i_i_o2_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNIMPSBK_LC_9_3_1 .C_ON=1'b0;
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNIMPSBK_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_10_c_RNIMPSBK_LC_9_3_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \sb_translator_1.state56_a_5_cry_10_c_RNIMPSBK_LC_9_3_1  (
            .in0(N__22450),
            .in1(N__22444),
            .in2(N__22438),
            .in3(N__22435),
            .lcout(),
            .ltout(\sb_translator_1.N_318_i_i_o2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_RNI41J131_7_LC_9_3_2 .C_ON=1'b0;
    defparam \sb_translator_1.state_RNI41J131_7_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_RNI41J131_7_LC_9_3_2 .LUT_INIT=16'b1011101110110011;
    LogicCell40 \sb_translator_1.state_RNI41J131_7_LC_9_3_2  (
            .in0(N__22151),
            .in1(N__22426),
            .in2(N__22369),
            .in3(N__22834),
            .lcout(\sb_translator_1.N_712 ),
            .ltout(\sb_translator_1.N_712_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_7_LC_9_3_3 .C_ON=1'b0;
    defparam \sb_translator_1.state_7_LC_9_3_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.state_7_LC_9_3_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \sb_translator_1.state_7_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22366),
            .in3(N__22347),
            .lcout(\sb_translator_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27461),
            .ce(),
            .sr(N__27087));
    defparam \sb_translator_1.cnt_leds_RNI8VOI7_0_LC_9_3_4 .C_ON=1'b0;
    defparam \sb_translator_1.cnt_leds_RNI8VOI7_0_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.cnt_leds_RNI8VOI7_0_LC_9_3_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \sb_translator_1.cnt_leds_RNI8VOI7_0_LC_9_3_4  (
            .in0(N__22135),
            .in1(N__22129),
            .in2(N__22123),
            .in3(N__22111),
            .lcout(\sb_translator_1.N_318_i_i_o2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_0_LC_9_3_5 .C_ON=1'b0;
    defparam \sb_translator_1.state_0_LC_9_3_5 .SEQ_MODE=4'b1011;
    defparam \sb_translator_1.state_0_LC_9_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \sb_translator_1.state_0_LC_9_3_5  (
            .in0(N__22099),
            .in1(N__21856),
            .in2(N__22828),
            .in3(N__22081),
            .lcout(\sb_translator_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27461),
            .ce(),
            .sr(N__27087));
    defparam \sb_translator_1.state_6_LC_9_4_0 .C_ON=1'b0;
    defparam \sb_translator_1.state_6_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.state_6_LC_9_4_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \sb_translator_1.state_6_LC_9_4_0  (
            .in0(N__22821),
            .in1(N__22752),
            .in2(N__22645),
            .in3(N__21855),
            .lcout(\sb_translator_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27470),
            .ce(),
            .sr(N__27093));
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNICLCM7_LC_9_4_1 .C_ON=1'b0;
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNICLCM7_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_13_c_RNICLCM7_LC_9_4_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \sb_translator_1.state56_a_5_cry_13_c_RNICLCM7_LC_9_4_1  (
            .in0(N__21835),
            .in1(N__21829),
            .in2(N__21823),
            .in3(N__21814),
            .lcout(),
            .ltout(\sb_translator_1.N_318_i_i_o2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIINPVD_LC_9_4_2 .C_ON=1'b0;
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIINPVD_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state56_a_5_cry_12_c_RNIINPVD_LC_9_4_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \sb_translator_1.state56_a_5_cry_12_c_RNIINPVD_LC_9_4_2  (
            .in0(N__22855),
            .in1(N__22849),
            .in2(N__22843),
            .in3(N__22840),
            .lcout(\sb_translator_1.N_318_i_i_o2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.state_1_LC_9_4_3 .C_ON=1'b0;
    defparam \sb_translator_1.state_1_LC_9_4_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.state_1_LC_9_4_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \sb_translator_1.state_1_LC_9_4_3  (
            .in0(N__22639),
            .in1(_gnd_net_),
            .in2(N__22784),
            .in3(N__22820),
            .lcout(\sb_translator_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27470),
            .ce(),
            .sr(N__27093));
    defparam \sb_translator_1.state_ns_i_i_0_0_o3_0_LC_9_4_4 .C_ON=1'b0;
    defparam \sb_translator_1.state_ns_i_i_0_0_o3_0_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.state_ns_i_i_0_0_o3_0_LC_9_4_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \sb_translator_1.state_ns_i_i_0_0_o3_0_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__22751),
            .in2(_gnd_net_),
            .in3(N__22638),
            .lcout(\sb_translator_1.state_ns_i_i_0_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_3_LC_9_5_0 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_3_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \ws2812.rgb_counter_3_LC_9_5_0 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \ws2812.rgb_counter_3_LC_9_5_0  (
            .in0(N__27750),
            .in1(N__27864),
            .in2(N__27607),
            .in3(N__26473),
            .lcout(\ws2812.rgb_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27476),
            .ce(),
            .sr(N__27098));
    defparam \ws2812.rgb_counter_0_LC_9_5_1 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_LC_9_5_1 .SEQ_MODE=4'b1011;
    defparam \ws2812.rgb_counter_0_LC_9_5_1 .LUT_INIT=16'b1110111000010001;
    LogicCell40 \ws2812.rgb_counter_0_LC_9_5_1  (
            .in0(N__27862),
            .in1(N__27749),
            .in2(_gnd_net_),
            .in3(N__27911),
            .lcout(\ws2812.rgb_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27476),
            .ce(),
            .sr(N__27098));
    defparam \ws2812.bit_counter_0_1_LC_9_5_2 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_1_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_0_1_LC_9_5_2 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \ws2812.bit_counter_0_1_LC_9_5_2  (
            .in0(N__27574),
            .in1(N__27863),
            .in2(_gnd_net_),
            .in3(N__24721),
            .lcout(\ws2812.bit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27476),
            .ce(),
            .sr(N__27098));
    defparam \sb_translator_1.addr_out_RNO_0_4_LC_9_5_4 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_4_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_4_LC_9_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_4_LC_9_5_4  (
            .in0(N__22582),
            .in1(N__22978),
            .in2(_gnd_net_),
            .in3(N__22564),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_RNO_0_6_LC_9_5_6 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_6_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_6_LC_9_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_6_LC_9_5_6  (
            .in0(N__22525),
            .in1(N__22507),
            .in2(_gnd_net_),
            .in3(N__22979),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.addr_out_RNO_0_7_LC_9_5_7 .C_ON=1'b0;
    defparam \sb_translator_1.addr_out_RNO_0_7_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \sb_translator_1.addr_out_RNO_0_7_LC_9_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \sb_translator_1.addr_out_RNO_0_7_LC_9_5_7  (
            .in0(N__22980),
            .in1(N__22944),
            .in2(_gnd_net_),
            .in3(N__22926),
            .lcout(\sb_translator_1.addr_out_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNING643_4_LC_9_6_0 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNING643_4_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNING643_4_LC_9_6_0 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \ws2812.bit_counter_0_RNING643_4_LC_9_6_0  (
            .in0(N__25400),
            .in1(N__26407),
            .in2(N__27747),
            .in3(N__26898),
            .lcout(\ws2812.bit_counter_0_RNING643Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNO_0_5_LC_9_6_1 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNO_0_5_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNO_0_5_LC_9_6_1 .LUT_INIT=16'b0111100001011010;
    LogicCell40 \ws2812.bit_counter_0_RNO_0_5_LC_9_6_1  (
            .in0(N__26899),
            .in1(N__27723),
            .in2(N__25231),
            .in3(N__25401),
            .lcout(\ws2812.un1_bit_counter_12_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNI6OQB3_2_LC_9_6_2 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNI6OQB3_2_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNI6OQB3_2_LC_9_6_2 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \ws2812.bit_counter_RNI6OQB3_2_LC_9_6_2  (
            .in0(N__25396),
            .in1(N__24664),
            .in2(N__27745),
            .in3(N__26894),
            .lcout(\ws2812.bit_counter_RNI6OQB3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNI7PQB3_3_LC_9_6_3 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNI7PQB3_3_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNI7PQB3_3_LC_9_6_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \ws2812.bit_counter_RNI7PQB3_3_LC_9_6_3  (
            .in0(N__26895),
            .in1(N__27715),
            .in2(N__24619),
            .in3(N__25397),
            .lcout(\ws2812.bit_counter_RNI7PQB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNI8QQB3_4_LC_9_6_4 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNI8QQB3_4_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNI8QQB3_4_LC_9_6_4 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \ws2812.bit_counter_RNI8QQB3_4_LC_9_6_4  (
            .in0(N__25399),
            .in1(N__24838),
            .in2(N__27746),
            .in3(N__26896),
            .lcout(\ws2812.bit_counter_RNI8QQB3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNI9RQB3_5_LC_9_6_5 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNI9RQB3_5_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNI9RQB3_5_LC_9_6_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \ws2812.bit_counter_RNI9RQB3_5_LC_9_6_5  (
            .in0(N__26897),
            .in1(N__27719),
            .in2(N__26368),
            .in3(N__25398),
            .lcout(\ws2812.bit_counter_RNI9RQB3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.new_data_req_RNO_0_LC_9_6_6 .C_ON=1'b0;
    defparam \ws2812.new_data_req_RNO_0_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.new_data_req_RNO_0_LC_9_6_6 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \ws2812.new_data_req_RNO_0_LC_9_6_6  (
            .in0(N__25402),
            .in1(N__27600),
            .in2(N__27748),
            .in3(N__26900),
            .lcout(),
            .ltout(\ws2812.N_140_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.new_data_req_LC_9_6_7 .C_ON=1'b0;
    defparam \ws2812.new_data_req_LC_9_6_7 .SEQ_MODE=4'b1010;
    defparam \ws2812.new_data_req_LC_9_6_7 .LUT_INIT=16'b1111111010101100;
    LogicCell40 \ws2812.new_data_req_LC_9_6_7  (
            .in0(N__22888),
            .in1(N__22869),
            .in2(N__22876),
            .in3(N__25403),
            .lcout(ws2812_next_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27484),
            .ce(),
            .sr(N__27103));
    defparam \sb_translator_1.rgb_data_out_0_LC_9_7_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_0_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_0_LC_9_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_0_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23182),
            .lcout(rgb_data_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \sb_translator_1.rgb_data_out_10_LC_9_7_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_10_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_10_LC_9_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.rgb_data_out_10_LC_9_7_1  (
            .in0(N__23173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_data_out_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \sb_translator_1.rgb_data_out_12_LC_9_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_12_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_12_LC_9_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_12_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23164),
            .lcout(rgb_data_out_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \sb_translator_1.rgb_data_out_18_LC_9_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_18_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_18_LC_9_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_18_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23155),
            .lcout(rgb_data_out_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \sb_translator_1.rgb_data_out_15_LC_9_7_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_15_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_15_LC_9_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_15_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23146),
            .lcout(rgb_data_out_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \sb_translator_1.rgb_data_out_16_LC_9_7_7 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_16_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_16_LC_9_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_16_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(rgb_data_out_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27490),
            .ce(N__27193),
            .sr(N__27111));
    defparam \demux.N_418_i_0_o2_0_LC_9_8_0 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_0_LC_9_8_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_418_i_0_o2_0_LC_9_8_0  (
            .in0(N__23125),
            .in1(N__23365),
            .in2(N__23434),
            .in3(N__23116),
            .lcout(),
            .ltout(\demux.N_418_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_1_LC_9_8_1 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_1_LC_9_8_1 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \demux.N_418_i_0_o2_1_LC_9_8_1  (
            .in0(N__23488),
            .in1(_gnd_net_),
            .in2(N__23110),
            .in3(N__23107),
            .lcout(),
            .ltout(\demux.N_418_i_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_o2_7_LC_9_8_2 .C_ON=1'b0;
    defparam \demux.N_418_i_0_o2_7_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_o2_7_LC_9_8_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \demux.N_418_i_0_o2_7_LC_9_8_2  (
            .in0(N__23089),
            .in1(N__23512),
            .in2(N__23077),
            .in3(N__23071),
            .lcout(\demux.N_418_i_0_o2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_418_i_0_a3_5_LC_9_8_3 .C_ON=1'b0;
    defparam \demux.N_418_i_0_a3_5_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_a3_5_LC_9_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_418_i_0_a3_5_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__23524),
            .in2(_gnd_net_),
            .in3(N__23293),
            .lcout(\demux.N_880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_0_LC_9_8_4 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_0_LC_9_8_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_420_i_0_o2_0_LC_9_8_4  (
            .in0(N__23506),
            .in1(N__23487),
            .in2(N__23433),
            .in3(N__23377),
            .lcout(),
            .ltout(\demux.N_420_i_0_o2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_1_LC_9_8_5 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_1_LC_9_8_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \demux.N_420_i_0_o2_1_LC_9_8_5  (
            .in0(N__23366),
            .in1(_gnd_net_),
            .in2(N__23317),
            .in3(N__23314),
            .lcout(),
            .ltout(\demux.N_420_i_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_7_LC_9_8_6 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_7_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_7_LC_9_8_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_420_i_0_o2_7_LC_9_8_6  (
            .in0(N__23294),
            .in1(N__23236),
            .in2(N__23221),
            .in3(N__23218),
            .lcout(\demux.N_420_i_0_o2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_a3_LC_9_9_1 .C_ON=1'b0;
    defparam \demux.N_417_i_0_a3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_a3_LC_9_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_417_i_0_a3_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__23209),
            .in2(_gnd_net_),
            .in3(N__25854),
            .lcout(\demux.N_888 ),
            .ltout(\demux.N_888_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_7_LC_9_9_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_7_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_7_LC_9_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_7_LC_9_9_2  (
            .in0(N__23883),
            .in1(N__23779),
            .in2(N__23197),
            .in3(N__23699),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27502),
            .ce(N__25437),
            .sr(N__27127));
    defparam \sb_translator_1.rgb_data_tmp_3_LC_9_9_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_3_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_3_LC_9_9_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_3_LC_9_9_3  (
            .in0(N__25859),
            .in1(N__24256),
            .in2(N__24218),
            .in3(N__24172),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27502),
            .ce(N__25437),
            .sr(N__27127));
    defparam \sb_translator_1.rgb_data_tmp_1_LC_9_9_4 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_1_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_1_LC_9_9_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_1_LC_9_9_4  (
            .in0(N__25855),
            .in1(N__24131),
            .in2(N__24085),
            .in3(N__24046),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27502),
            .ce(N__25437),
            .sr(N__27127));
    defparam \demux.N_418_i_0_a3_LC_9_9_5 .C_ON=1'b0;
    defparam \demux.N_418_i_0_a3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_418_i_0_a3_LC_9_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_418_i_0_a3_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__23194),
            .in2(_gnd_net_),
            .in3(N__25852),
            .lcout(\demux.N_874 ),
            .ltout(\demux.N_874_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_6_LC_9_9_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_6_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_6_LC_9_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_6_LC_9_9_6  (
            .in0(N__23618),
            .in1(N__23582),
            .in2(N__23797),
            .in3(N__23551),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27502),
            .ce(N__25437),
            .sr(N__27127));
    defparam \demux.N_420_i_0_a3_LC_9_9_7 .C_ON=1'b0;
    defparam \demux.N_420_i_0_a3_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_a3_LC_9_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_420_i_0_a3_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__23794),
            .in2(_gnd_net_),
            .in3(N__25853),
            .lcout(\demux.N_420_i_0_aZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_tmp_23_LC_9_10_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_23_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_23_LC_9_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_23_LC_9_10_0  (
            .in0(N__23721),
            .in1(N__23882),
            .in2(N__23701),
            .in3(N__23770),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27507),
            .ce(N__25077),
            .sr(N__27130));
    defparam \sb_translator_1.rgb_data_tmp_22_LC_9_10_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_22_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_22_LC_9_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_22_LC_9_10_1  (
            .in0(N__23625),
            .in1(N__23595),
            .in2(N__23658),
            .in3(N__23559),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27507),
            .ce(N__25077),
            .sr(N__27130));
    defparam \sb_translator_1.rgb_data_tmp_21_LC_9_10_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_21_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_21_LC_9_10_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_21_LC_9_10_2  (
            .in0(N__25850),
            .in1(N__25757),
            .in2(N__25715),
            .in3(N__25656),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27507),
            .ce(N__25077),
            .sr(N__27130));
    defparam \sb_translator_1.rgb_data_tmp_19_LC_9_10_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_19_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_19_LC_9_10_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_19_LC_9_10_3  (
            .in0(N__24211),
            .in1(N__24264),
            .in2(N__25867),
            .in3(N__24176),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27507),
            .ce(N__25077),
            .sr(N__27130));
    defparam \sb_translator_1.rgb_data_tmp_17_LC_9_10_5 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_17_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_17_LC_9_10_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \sb_translator_1.rgb_data_tmp_17_LC_9_10_5  (
            .in0(N__24093),
            .in1(N__25851),
            .in2(N__24136),
            .in3(N__24043),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27507),
            .ce(N__25077),
            .sr(N__27130));
    defparam \sb_translator_1.instr_out_7_LC_9_11_0 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_7_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_7_LC_9_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.instr_out_7_LC_9_11_0  (
            .in0(N__23881),
            .in1(N__23778),
            .in2(N__23725),
            .in3(N__23698),
            .lcout(miso_data_in_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \sb_translator_1.instr_out_6_LC_9_11_1 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_6_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_6_LC_9_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.instr_out_6_LC_9_11_1  (
            .in0(N__23659),
            .in1(N__23629),
            .in2(N__23599),
            .in3(N__23560),
            .lcout(miso_data_in_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \sb_translator_1.instr_out_5_LC_9_11_2 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_5_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_5_LC_9_11_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.instr_out_5_LC_9_11_2  (
            .in0(N__25861),
            .in1(N__25765),
            .in2(N__25711),
            .in3(N__25654),
            .lcout(miso_data_in_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \sb_translator_1.instr_out_3_LC_9_11_3 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_3_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_3_LC_9_11_3 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \sb_translator_1.instr_out_3_LC_9_11_3  (
            .in0(N__24265),
            .in1(N__24219),
            .in2(N__24178),
            .in3(N__25862),
            .lcout(miso_data_in_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \sb_translator_1.instr_out_1_LC_9_11_4 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_1_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_1_LC_9_11_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.instr_out_1_LC_9_11_4  (
            .in0(N__25860),
            .in1(N__24135),
            .in2(N__24097),
            .in3(N__24045),
            .lcout(miso_data_in_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \sb_translator_1.instr_out_4_LC_9_11_5 .C_ON=1'b0;
    defparam \sb_translator_1.instr_out_4_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.instr_out_4_LC_9_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.instr_out_4_LC_9_11_5  (
            .in0(N__25603),
            .in1(N__25581),
            .in2(N__25540),
            .in3(N__25484),
            .lcout(miso_data_in_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27511),
            .ce(N__23991),
            .sr(N__27134));
    defparam \demux.N_417_i_0_a3_7_LC_9_12_0 .C_ON=1'b0;
    defparam \demux.N_417_i_0_a3_7_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_a3_7_LC_9_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \demux.N_417_i_0_a3_7_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__23971),
            .in2(_gnd_net_),
            .in3(N__23955),
            .lcout(),
            .ltout(\demux.N_417_i_0_a3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_8_LC_9_12_1 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_8_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_8_LC_9_12_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \demux.N_417_i_0_o2_8_LC_9_12_1  (
            .in0(N__23899),
            .in1(N__23839),
            .in2(N__23887),
            .in3(N__24358),
            .lcout(\demux.N_417_i_0_o2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_417_i_0_o2_4_LC_9_12_3 .C_ON=1'b0;
    defparam \demux.N_417_i_0_o2_4_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \demux.N_417_i_0_o2_4_LC_9_12_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_417_i_0_o2_4_LC_9_12_3  (
            .in0(N__24432),
            .in1(N__23857),
            .in2(N__24508),
            .in3(N__23845),
            .lcout(\demux.N_417_i_0_o2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_422_i_0_o2_4_LC_9_12_4 .C_ON=1'b0;
    defparam \demux.N_422_i_0_o2_4_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \demux.N_422_i_0_o2_4_LC_9_12_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_422_i_0_o2_4_LC_9_12_4  (
            .in0(N__23833),
            .in1(N__24502),
            .in2(N__23824),
            .in3(N__24431),
            .lcout(\demux.N_422_i_0_o2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_419_i_0_o2_4_LC_9_12_5 .C_ON=1'b0;
    defparam \demux.N_419_i_0_o2_4_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \demux.N_419_i_0_o2_4_LC_9_12_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \demux.N_419_i_0_o2_4_LC_9_12_5  (
            .in0(N__24430),
            .in1(N__24544),
            .in2(N__24507),
            .in3(N__24532),
            .lcout(\demux.N_419_i_0_o2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_4_LC_9_12_6 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_4_LC_9_12_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \demux.N_420_i_0_o2_4_LC_9_12_6  (
            .in0(N__24520),
            .in1(N__24503),
            .in2(N__24451),
            .in3(N__24433),
            .lcout(),
            .ltout(\demux.N_420_i_0_o2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \demux.N_420_i_0_o2_8_LC_9_12_7 .C_ON=1'b0;
    defparam \demux.N_420_i_0_o2_8_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \demux.N_420_i_0_o2_8_LC_9_12_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \demux.N_420_i_0_o2_8_LC_9_12_7  (
            .in0(N__24376),
            .in1(N__24359),
            .in2(N__24292),
            .in3(N__24289),
            .lcout(\demux.N_420_i_0_o2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIKD643_1_LC_11_3_0 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIKD643_1_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIKD643_1_LC_11_3_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \ws2812.bit_counter_0_RNIKD643_1_LC_11_3_0  (
            .in0(N__27734),
            .in1(N__26860),
            .in2(N__24769),
            .in3(N__25360),
            .lcout(\ws2812.bit_counter_0_RNIKD643Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNILE643_2_LC_11_3_1 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNILE643_2_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNILE643_2_LC_11_3_1 .LUT_INIT=16'b1010101000001010;
    LogicCell40 \ws2812.bit_counter_0_RNILE643_2_LC_11_3_1  (
            .in0(N__26861),
            .in1(N__24895),
            .in2(N__25393),
            .in3(N__27735),
            .lcout(\ws2812.bit_counter_0_RNILE643Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIMF643_3_LC_11_3_2 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIMF643_3_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIMF643_3_LC_11_3_2 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ws2812.bit_counter_0_RNIMF643_3_LC_11_3_2  (
            .in0(N__27736),
            .in1(N__25361),
            .in2(N__24868),
            .in3(N__26862),
            .lcout(\ws2812.bit_counter_0_RNIMF643Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.state_1_LC_11_3_3 .C_ON=1'b0;
    defparam \ws2812.state_1_LC_11_3_3 .SEQ_MODE=4'b1010;
    defparam \ws2812.state_1_LC_11_3_3 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \ws2812.state_1_LC_11_3_3  (
            .in0(N__26863),
            .in1(N__27786),
            .in2(N__25394),
            .in3(N__27737),
            .lcout(\ws2812.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27471),
            .ce(),
            .sr(N__27094));
    defparam \ws2812.un1_bit_counter_12_cry_0_c_RNO_LC_11_3_4 .C_ON=1'b0;
    defparam \ws2812.un1_bit_counter_12_cry_0_c_RNO_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.un1_bit_counter_12_cry_0_c_RNO_LC_11_3_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ws2812.un1_bit_counter_12_cry_0_c_RNO_LC_11_3_4  (
            .in0(N__27732),
            .in1(N__25355),
            .in2(N__25275),
            .in3(N__26858),
            .lcout(\ws2812.un1_bit_counter_12_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNI5NQB3_1_LC_11_3_6 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNI5NQB3_1_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNI5NQB3_1_LC_11_3_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \ws2812.bit_counter_RNI5NQB3_1_LC_11_3_6  (
            .in0(N__27733),
            .in1(N__26859),
            .in2(N__25303),
            .in3(N__25356),
            .lcout(\ws2812.bit_counter_RNI5NQB3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNIENHA_3_LC_11_4_0 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNIENHA_3_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNIENHA_3_LC_11_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_RNIENHA_3_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24607),
            .lcout(\ws2812.un6_data_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIQAT2_0_LC_11_4_1 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIQAT2_0_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIQAT2_0_LC_11_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_0_RNIQAT2_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25181),
            .lcout(\ws2812.bit_counter_0_RNIQAT2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIRBT2_1_LC_11_4_2 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIRBT2_1_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIRBT2_1_LC_11_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_0_RNIRBT2_1_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24765),
            .lcout(\ws2812.bit_counter_0_RNIRBT2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIG4UQ_0_LC_11_4_3 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIG4UQ_0_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIG4UQ_0_LC_11_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ws2812.bit_counter_0_RNIG4UQ_0_LC_11_4_3  (
            .in0(N__24764),
            .in1(N__24655),
            .in2(N__24612),
            .in3(N__25180),
            .lcout(\ws2812.state_ns_0_i_o2_6_0 ),
            .ltout(\ws2812.state_ns_0_i_o2_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNISPQG2_0_LC_11_4_4 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNISPQG2_0_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNISPQG2_0_LC_11_4_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ws2812.bit_counter_0_RNISPQG2_0_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__25311),
            .in2(N__24568),
            .in3(N__24906),
            .lcout(\ws2812.N_105 ),
            .ltout(\ws2812.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIJC643_0_LC_11_4_5 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIJC643_0_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIJC643_0_LC_11_4_5 .LUT_INIT=16'b1011000010110000;
    LogicCell40 \ws2812.bit_counter_0_RNIJC643_0_LC_11_4_5  (
            .in0(N__27741),
            .in1(N__25369),
            .in2(N__24565),
            .in3(N__25182),
            .lcout(\ws2812.bit_counter_0_RNIJC643Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.state_RNIBU1P2_1_LC_11_4_6 .C_ON=1'b0;
    defparam \ws2812.state_RNIBU1P2_1_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.state_RNIBU1P2_1_LC_11_4_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ws2812.state_RNIBU1P2_1_LC_11_4_6  (
            .in0(N__24562),
            .in1(N__25312),
            .in2(N__25395),
            .in3(N__24907),
            .lcout(\ws2812.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNIDMHA_2_LC_11_4_7 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNIDMHA_2_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNIDMHA_2_LC_11_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_RNIDMHA_2_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24656),
            .lcout(\ws2812.un6_data_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un1_bit_counter_12_cry_0_c_LC_11_5_0 .C_ON=1'b1;
    defparam \ws2812.un1_bit_counter_12_cry_0_c_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.un1_bit_counter_12_cry_0_c_LC_11_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ws2812.un1_bit_counter_12_cry_0_c_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__25270),
            .in2(N__24556),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\ws2812.un1_bit_counter_12_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_1_LC_11_5_1 .C_ON=1'b1;
    defparam \ws2812.bit_counter_1_LC_11_5_1 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_1_LC_11_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_1_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__25296),
            .in2(N__24793),
            .in3(N__24781),
            .lcout(\ws2812.bit_counterZ0Z_1 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_0 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_1 ),
            .clk(N__27485),
            .ce(),
            .sr(N__27108));
    defparam \ws2812.bit_counter_0_RNO_0_0_LC_11_5_2 .C_ON=1'b1;
    defparam \ws2812.bit_counter_0_RNO_0_0_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNO_0_0_LC_11_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_0_RNO_0_0_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__24778),
            .in2(N__25189),
            .in3(N__24772),
            .lcout(\ws2812.bit_counter_0_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_1 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNO_0_1_LC_11_5_3 .C_ON=1'b1;
    defparam \ws2812.bit_counter_0_RNO_0_1_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNO_0_1_LC_11_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_0_RNO_0_1_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__24760),
            .in2(N__24733),
            .in3(N__24712),
            .lcout(\ws2812.bit_counter_0_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_2 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_2_LC_11_5_4 .C_ON=1'b1;
    defparam \ws2812.bit_counter_0_2_LC_11_5_4 .SEQ_MODE=4'b1011;
    defparam \ws2812.bit_counter_0_2_LC_11_5_4 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \ws2812.bit_counter_0_2_LC_11_5_4  (
            .in0(N__27828),
            .in1(N__24889),
            .in2(N__24709),
            .in3(N__24697),
            .lcout(\ws2812.bit_counterZ0Z_4 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_3 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_4 ),
            .clk(N__27485),
            .ce(),
            .sr(N__27108));
    defparam \ws2812.bit_counter_0_3_LC_11_5_5 .C_ON=1'b1;
    defparam \ws2812.bit_counter_0_3_LC_11_5_5 .SEQ_MODE=4'b1011;
    defparam \ws2812.bit_counter_0_3_LC_11_5_5 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \ws2812.bit_counter_0_3_LC_11_5_5  (
            .in0(N__27855),
            .in1(N__24859),
            .in2(N__24694),
            .in3(N__24682),
            .lcout(\ws2812.bit_counterZ0Z_5 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_4 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_5 ),
            .clk(N__27485),
            .ce(),
            .sr(N__27108));
    defparam \ws2812.bit_counter_2_LC_11_5_6 .C_ON=1'b1;
    defparam \ws2812.bit_counter_2_LC_11_5_6 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_2_LC_11_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_2_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__24657),
            .in2(N__24679),
            .in3(N__24637),
            .lcout(\ws2812.bit_counter_6 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_5 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_6 ),
            .clk(N__27485),
            .ce(),
            .sr(N__27108));
    defparam \ws2812.bit_counter_3_LC_11_5_7 .C_ON=1'b1;
    defparam \ws2812.bit_counter_3_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_3_LC_11_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_3_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__24608),
            .in2(N__24634),
            .in3(N__24586),
            .lcout(\ws2812.bit_counter_7 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_6 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_7 ),
            .clk(N__27485),
            .ce(),
            .sr(N__27108));
    defparam \ws2812.bit_counter_4_LC_11_6_0 .C_ON=1'b1;
    defparam \ws2812.bit_counter_4_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_4_LC_11_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_4_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__24834),
            .in2(N__24583),
            .in3(N__24571),
            .lcout(\ws2812.bit_counter_8 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\ws2812.un1_bit_counter_12_cry_8 ),
            .clk(N__27493),
            .ce(),
            .sr(N__27112));
    defparam \ws2812.bit_counter_5_LC_11_6_1 .C_ON=1'b1;
    defparam \ws2812.bit_counter_5_LC_11_6_1 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_5_LC_11_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_5_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__26354),
            .in2(N__24949),
            .in3(N__24937),
            .lcout(\ws2812.bit_counter_9 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_8 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_9 ),
            .clk(N__27493),
            .ce(),
            .sr(N__27112));
    defparam \ws2812.bit_counter_0_RNO_0_4_LC_11_6_2 .C_ON=1'b1;
    defparam \ws2812.bit_counter_0_RNO_0_4_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNO_0_4_LC_11_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.bit_counter_0_RNO_0_4_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__26403),
            .in2(N__24934),
            .in3(N__24922),
            .lcout(\ws2812.bit_counter_0_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\ws2812.un1_bit_counter_12_cry_9 ),
            .carryout(\ws2812.un1_bit_counter_12_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_5_LC_11_6_3 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_5_LC_11_6_3 .SEQ_MODE=4'b1011;
    defparam \ws2812.bit_counter_0_5_LC_11_6_3 .LUT_INIT=16'b1011101011101010;
    LogicCell40 \ws2812.bit_counter_0_5_LC_11_6_3  (
            .in0(N__27575),
            .in1(N__24919),
            .in2(N__27865),
            .in3(N__24910),
            .lcout(\ws2812.bit_counter_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27493),
            .ce(),
            .sr(N__27112));
    defparam \ws2812.bit_counter_0_RNIOCUQ_2_LC_11_7_0 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIOCUQ_2_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIOCUQ_2_LC_11_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ws2812.bit_counter_0_RNIOCUQ_2_LC_11_7_0  (
            .in0(N__24893),
            .in1(N__24832),
            .in2(N__26364),
            .in3(N__24863),
            .lcout(\ws2812.state_ns_0_i_o2_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNISCT2_2_LC_11_7_1 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNISCT2_2_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNISCT2_2_LC_11_7_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ws2812.bit_counter_0_RNISCT2_2_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__24894),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ws2812.bit_counter_0_RNISCT2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNITDT2_3_LC_11_7_2 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNITDT2_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNITDT2_3_LC_11_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_0_RNITDT2_3_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24864),
            .lcout(\ws2812.bit_counter_0_RNITDT2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNIFOHA_4_LC_11_7_3 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNIFOHA_4_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNIFOHA_4_LC_11_7_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ws2812.bit_counter_RNIFOHA_4_LC_11_7_3  (
            .in0(N__24833),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ws2812.un6_data_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_0_LC_11_7_5 .C_ON=1'b0;
    defparam \ws2812.data_RNO_0_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_0_LC_11_7_5 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \ws2812.data_RNO_0_LC_11_7_5  (
            .in0(N__26242),
            .in1(N__24982),
            .in2(N__25906),
            .in3(N__26542),
            .lcout(),
            .ltout(\ws2812.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_LC_11_7_6 .C_ON=1'b0;
    defparam \ws2812.data_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \ws2812.data_LC_11_7_6 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \ws2812.data_LC_11_7_6  (
            .in0(N__24804),
            .in1(N__25407),
            .in2(N__24814),
            .in3(N__26296),
            .lcout(led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27498),
            .ce(),
            .sr(N__27123));
    defparam \ws2812.data_RNO_7_LC_11_7_7 .C_ON=1'b0;
    defparam \ws2812.data_RNO_7_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_7_LC_11_7_7 .LUT_INIT=16'b0101011100000011;
    LogicCell40 \ws2812.data_RNO_7_LC_11_7_7  (
            .in0(N__26241),
            .in1(N__25276),
            .in2(N__25905),
            .in3(N__24981),
            .lcout(\ws2812.N_135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI2H7O_2_LC_11_8_0 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI2H7O_2_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI2H7O_2_LC_11_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ws2812.rgb_counter_RNI2H7O_2_LC_11_8_0  (
            .in0(N__25039),
            .in1(N__24955),
            .in2(_gnd_net_),
            .in3(N__28114),
            .lcout(\ws2812.rgb_counter_RNI2H7OZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIFI3M_2_LC_11_8_1 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIFI3M_2_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIFI3M_2_LC_11_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ws2812.rgb_counter_RNIFI3M_2_LC_11_8_1  (
            .in0(N__28115),
            .in1(N__25027),
            .in2(_gnd_net_),
            .in3(N__25135),
            .lcout(\ws2812.rgb_counter_RNIFI3MZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIDG3M_2_LC_11_8_2 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIDG3M_2_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIDG3M_2_LC_11_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ws2812.rgb_counter_RNIDG3M_2_LC_11_8_2  (
            .in0(N__26587),
            .in1(N__25015),
            .in2(_gnd_net_),
            .in3(N__28117),
            .lcout(),
            .ltout(\ws2812.rgb_counter_RNIDG3MZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIUE972_1_LC_11_8_3 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIUE972_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIUE972_1_LC_11_8_3 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ws2812.rgb_counter_RNIUE972_1_LC_11_8_3  (
            .in0(N__28033),
            .in1(N__27933),
            .in2(N__25003),
            .in3(N__25000),
            .lcout(),
            .ltout(\ws2812.rgb_data_pmux_22_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIOQ324_0_LC_11_8_4 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIOQ324_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIOQ324_0_LC_11_8_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ws2812.rgb_counter_RNIOQ324_0_LC_11_8_4  (
            .in0(N__27934),
            .in1(N__24994),
            .in2(N__24988),
            .in3(N__24973),
            .lcout(),
            .ltout(\ws2812.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI0NBTB_3_LC_11_8_5 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI0NBTB_3_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI0NBTB_3_LC_11_8_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ws2812.rgb_counter_RNI0NBTB_3_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__27994),
            .in2(N__24985),
            .in3(N__26533),
            .lcout(\ws2812.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI4J7O_2_LC_11_8_6 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI4J7O_2_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI4J7O_2_LC_11_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ws2812.rgb_counter_RNI4J7O_2_LC_11_8_6  (
            .in0(N__25153),
            .in1(N__25114),
            .in2(_gnd_net_),
            .in3(N__28116),
            .lcout(\ws2812.rgb_counter_RNI4J7OZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_out_8_LC_11_8_7 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_8_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_8_LC_11_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_8_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24967),
            .lcout(rgb_data_out_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27505),
            .ce(N__27194),
            .sr(N__27128));
    defparam \sb_translator_1.rgb_data_out_13_LC_11_9_0 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_13_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_13_LC_11_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_13_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25165),
            .lcout(rgb_data_out_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_11_LC_11_9_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_11_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_11_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_11_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25147),
            .lcout(rgb_data_out_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_4_LC_11_9_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_4_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_4_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_4_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25450),
            .lcout(rgb_data_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_9_LC_11_9_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_9_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_9_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_9_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25126),
            .lcout(rgb_data_out_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_5_LC_11_9_4 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_5_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_5_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_5_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25633),
            .lcout(rgb_data_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_20_LC_11_9_5 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_20_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_20_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_20_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25084),
            .lcout(rgb_data_out_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_1_LC_11_9_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_1_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_1_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_1_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25105),
            .lcout(rgb_data_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_out_21_LC_11_9_7 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_21_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_21_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_21_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25096),
            .lcout(rgb_data_out_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27508),
            .ce(N__27191),
            .sr(N__27131));
    defparam \sb_translator_1.rgb_data_tmp_20_LC_11_10_6 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_20_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_20_LC_11_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_20_LC_11_10_6  (
            .in0(N__25624),
            .in1(N__25570),
            .in2(N__25534),
            .in3(N__25485),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27514),
            .ce(N__25078),
            .sr(N__27135));
    defparam \sb_translator_1.rgb_data_tmp_5_LC_11_11_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_5_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_5_LC_11_11_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \sb_translator_1.rgb_data_tmp_5_LC_11_11_1  (
            .in0(N__25866),
            .in1(N__25764),
            .in2(N__25722),
            .in3(N__25663),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27516),
            .ce(N__25441),
            .sr(N__27137));
    defparam \sb_translator_1.rgb_data_tmp_4_LC_11_11_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_tmp_4_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_tmp_4_LC_11_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \sb_translator_1.rgb_data_tmp_4_LC_11_11_3  (
            .in0(N__25622),
            .in1(N__25582),
            .in2(N__25538),
            .in3(N__25486),
            .lcout(\sb_translator_1.rgb_data_tmpZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27516),
            .ce(N__25441),
            .sr(N__27137));
    defparam \ws2812.bit_counter_0_LC_12_3_7 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_LC_12_3_7 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_0_LC_12_3_7 .LUT_INIT=16'b0011101111000100;
    LogicCell40 \ws2812.bit_counter_0_LC_12_3_7  (
            .in0(N__25365),
            .in1(N__26872),
            .in2(N__27751),
            .in3(N__25274),
            .lcout(\ws2812.bit_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27479),
            .ce(),
            .sr(N__27099));
    defparam \ws2812.bit_counter_0_RNIK8UQ_5_LC_12_4_0 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIK8UQ_5_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIK8UQ_5_LC_12_4_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ws2812.bit_counter_0_RNIK8UQ_5_LC_12_4_0  (
            .in0(N__25294),
            .in1(N__26392),
            .in2(N__25230),
            .in3(N__25256),
            .lcout(\ws2812.state_ns_0_i_o2_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNICLHA_1_LC_12_4_1 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNICLHA_1_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNICLHA_1_LC_12_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_RNICLHA_1_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25295),
            .lcout(\ws2812.un6_data_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un6_data_cry_0_c_inv_LC_12_4_4 .C_ON=1'b0;
    defparam \ws2812.un6_data_cry_0_c_inv_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.un6_data_cry_0_c_inv_LC_12_4_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ws2812.un6_data_cry_0_c_inv_LC_12_4_4  (
            .in0(N__26171),
            .in1(N__25257),
            .in2(_gnd_net_),
            .in3(N__26290),
            .lcout(\ws2812.bit_counter_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIVFT2_5_LC_12_4_5 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIVFT2_5_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIVFT2_5_LC_12_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_0_RNIVFT2_5_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25226),
            .lcout(\ws2812.un6_data_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_4_LC_12_4_6 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_4_LC_12_4_6 .SEQ_MODE=4'b1011;
    defparam \ws2812.bit_counter_0_4_LC_12_4_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \ws2812.bit_counter_0_4_LC_12_4_6  (
            .in0(N__27829),
            .in1(N__27577),
            .in2(_gnd_net_),
            .in3(N__25204),
            .lcout(\ws2812.bit_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27486),
            .ce(),
            .sr(N__27109));
    defparam \ws2812.bit_counter_0_0_LC_12_4_7 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_0_LC_12_4_7 .SEQ_MODE=4'b1010;
    defparam \ws2812.bit_counter_0_0_LC_12_4_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \ws2812.bit_counter_0_0_LC_12_4_7  (
            .in0(N__27576),
            .in1(N__25195),
            .in2(_gnd_net_),
            .in3(N__27830),
            .lcout(\ws2812.bit_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27486),
            .ce(),
            .sr(N__27109));
    defparam \ws2812.un6_data_cry_0_c_LC_12_5_0 .C_ON=1'b1;
    defparam \ws2812.un6_data_cry_0_c_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.un6_data_cry_0_c_LC_12_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ws2812.un6_data_cry_0_c_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__26289),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\ws2812.un6_data_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_8_LC_12_5_1 .C_ON=1'b1;
    defparam \ws2812.data_RNO_8_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_8_LC_12_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_8_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__26278),
            .in2(_gnd_net_),
            .in3(N__26272),
            .lcout(\ws2812.data_RNOZ0Z_8 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_0 ),
            .carryout(\ws2812.un6_data_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_9_LC_12_5_2 .C_ON=1'b1;
    defparam \ws2812.data_RNO_9_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_9_LC_12_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.data_RNO_9_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__26269),
            .in2(N__26210),
            .in3(N__26263),
            .lcout(\ws2812.data_RNOZ0Z_9 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_1 ),
            .carryout(\ws2812.un6_data_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_10_LC_12_5_3 .C_ON=1'b1;
    defparam \ws2812.data_RNO_10_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_10_LC_12_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.data_RNO_10_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__26260),
            .in2(N__26208),
            .in3(N__26254),
            .lcout(\ws2812.data_RNOZ0Z_10 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_2 ),
            .carryout(\ws2812.un6_data_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un6_data_cry_3_c_RNIKNFB_LC_12_5_4 .C_ON=1'b1;
    defparam \ws2812.un6_data_cry_3_c_RNIKNFB_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.un6_data_cry_3_c_RNIKNFB_LC_12_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.un6_data_cry_3_c_RNIKNFB_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__26251),
            .in2(N__26211),
            .in3(N__26230),
            .lcout(\ws2812.un6_data_cry_3_c_RNIKNFBZ0 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_3 ),
            .carryout(\ws2812.un6_data_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un6_data_cry_4_c_RNIMQGB_LC_12_5_5 .C_ON=1'b1;
    defparam \ws2812.un6_data_cry_4_c_RNIMQGB_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.un6_data_cry_4_c_RNIMQGB_LC_12_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.un6_data_cry_4_c_RNIMQGB_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__26227),
            .in2(N__26209),
            .in3(N__25888),
            .lcout(\ws2812.un6_data_cry_4_c_RNIMQGBZ0 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_4 ),
            .carryout(\ws2812.un6_data_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_3_LC_12_5_6 .C_ON=1'b1;
    defparam \ws2812.data_RNO_3_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_3_LC_12_5_6 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \ws2812.data_RNO_3_LC_12_5_6  (
            .in0(N__27696),
            .in1(N__25885),
            .in2(_gnd_net_),
            .in3(N__25879),
            .lcout(\ws2812.data_5_iv_0_47_a2_0_a2_0 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_5 ),
            .carryout(\ws2812.un6_data_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_11_LC_12_5_7 .C_ON=1'b1;
    defparam \ws2812.data_RNO_11_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_11_LC_12_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_11_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__25876),
            .in2(_gnd_net_),
            .in3(N__25870),
            .lcout(\ws2812.data_RNOZ0Z_11 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_6 ),
            .carryout(\ws2812.un6_data_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_12_LC_12_6_0 .C_ON=1'b1;
    defparam \ws2812.data_RNO_12_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_12_LC_12_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_12_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__26458),
            .in2(_gnd_net_),
            .in3(N__26452),
            .lcout(\ws2812.data_RNOZ0Z_12 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\ws2812.un6_data_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_13_LC_12_6_1 .C_ON=1'b1;
    defparam \ws2812.data_RNO_13_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_13_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_13_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__26329),
            .in2(_gnd_net_),
            .in3(N__26449),
            .lcout(\ws2812.data_RNOZ0Z_13 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_8 ),
            .carryout(\ws2812.un6_data_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_5_LC_12_6_2 .C_ON=1'b1;
    defparam \ws2812.data_RNO_5_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_5_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_5_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__26374),
            .in2(_gnd_net_),
            .in3(N__26446),
            .lcout(\ws2812.data_RNOZ0Z_5 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_9 ),
            .carryout(\ws2812.un6_data_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_6_LC_12_6_3 .C_ON=1'b1;
    defparam \ws2812.data_RNO_6_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_6_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ws2812.data_RNO_6_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__26443),
            .in2(_gnd_net_),
            .in3(N__26434),
            .lcout(\ws2812.data_RNOZ0Z_6 ),
            .ltout(),
            .carryin(\ws2812.un6_data_cry_10 ),
            .carryout(\ws2812.un6_data_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_4_LC_12_6_4 .C_ON=1'b0;
    defparam \ws2812.data_RNO_4_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_4_LC_12_6_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ws2812.data_RNO_4_LC_12_6_4  (
            .in0(N__26431),
            .in1(N__26425),
            .in2(N__26419),
            .in3(N__26410),
            .lcout(\ws2812.data_5_iv_0_47_a2_0_a2_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_0_RNIUET2_4_LC_12_6_5 .C_ON=1'b0;
    defparam \ws2812.bit_counter_0_RNIUET2_4_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_0_RNIUET2_4_LC_12_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ws2812.bit_counter_0_RNIUET2_4_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\ws2812.un6_data_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.bit_counter_RNIGPHA_5_LC_12_6_6 .C_ON=1'b0;
    defparam \ws2812.bit_counter_RNIGPHA_5_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.bit_counter_RNIGPHA_5_LC_12_6_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \ws2812.bit_counter_RNIGPHA_5_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__26353),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ws2812.un6_data_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_1_LC_12_6_7 .C_ON=1'b0;
    defparam \ws2812.data_RNO_1_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_1_LC_12_6_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ws2812.data_RNO_1_LC_12_6_7  (
            .in0(N__26323),
            .in1(N__26317),
            .in2(N__26311),
            .in3(N__26302),
            .lcout(\ws2812.data_5_iv_0_47_a2_0_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.data_RNO_2_LC_12_7_1 .C_ON=1'b0;
    defparam \ws2812.data_RNO_2_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.data_RNO_2_LC_12_7_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ws2812.data_RNO_2_LC_12_7_1  (
            .in0(N__26578),
            .in1(N__26569),
            .in2(N__26560),
            .in3(N__26548),
            .lcout(\ws2812.data_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIVOJT3_1_LC_12_7_2 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIVOJT3_1_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIVOJT3_1_LC_12_7_2 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ws2812.rgb_counter_RNIVOJT3_1_LC_12_7_2  (
            .in0(N__28032),
            .in1(N__27931),
            .in2(N__26701),
            .in3(N__26485),
            .lcout(),
            .ltout(\ws2812.rgb_data_pmux_15_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIUIOE7_0_LC_12_7_3 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIUIOE7_0_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIUIOE7_0_LC_12_7_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ws2812.rgb_counter_RNIUIOE7_0_LC_12_7_3  (
            .in0(N__27932),
            .in1(N__26668),
            .in2(N__26536),
            .in3(N__26818),
            .lcout(\ws2812.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_0_RNIN42Q_3_LC_12_7_4 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_RNIN42Q_3_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_0_RNIN42Q_3_LC_12_7_4 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ws2812.rgb_counter_0_RNIN42Q_3_LC_12_7_4  (
            .in0(N__26754),
            .in1(N__28106),
            .in2(N__26527),
            .in3(N__26515),
            .lcout(),
            .ltout(\ws2812.rgb_data_pmux_3_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIKHAI1_2_LC_12_7_5 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIKHAI1_2_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIKHAI1_2_LC_12_7_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ws2812.rgb_counter_RNIKHAI1_2_LC_12_7_5  (
            .in0(N__28107),
            .in1(N__26506),
            .in2(N__26497),
            .in3(N__26494),
            .lcout(\ws2812.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un1_rgb_counter_cry_0_c_LC_12_8_0 .C_ON=1'b1;
    defparam \ws2812.un1_rgb_counter_cry_0_c_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.un1_rgb_counter_cry_0_c_LC_12_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ws2812.un1_rgb_counter_cry_0_c_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__27936),
            .in2(N__27874),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\ws2812.un1_rgb_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_1_LC_12_8_1 .C_ON=1'b1;
    defparam \ws2812.rgb_counter_1_LC_12_8_1 .SEQ_MODE=4'b1011;
    defparam \ws2812.rgb_counter_1_LC_12_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.rgb_counter_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__28035),
            .in2(N__28006),
            .in3(N__26479),
            .lcout(\ws2812.rgb_counterZ0Z_1 ),
            .ltout(),
            .carryin(\ws2812.un1_rgb_counter_cry_0 ),
            .carryout(\ws2812.un1_rgb_counter_cry_1 ),
            .clk(N__27509),
            .ce(),
            .sr(N__27132));
    defparam \ws2812.rgb_counter_2_LC_12_8_2 .C_ON=1'b1;
    defparam \ws2812.rgb_counter_2_LC_12_8_2 .SEQ_MODE=4'b1011;
    defparam \ws2812.rgb_counter_2_LC_12_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.rgb_counter_2_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__28118),
            .in2(N__28048),
            .in3(N__26476),
            .lcout(\ws2812.rgb_counterZ0Z_2 ),
            .ltout(),
            .carryin(\ws2812.un1_rgb_counter_cry_1 ),
            .carryout(\ws2812.un1_rgb_counter_cry_2 ),
            .clk(N__27509),
            .ce(),
            .sr(N__27132));
    defparam \ws2812.rgb_counter_RNO_0_3_LC_12_8_3 .C_ON=1'b1;
    defparam \ws2812.rgb_counter_RNO_0_3_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNO_0_3_LC_12_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ws2812.rgb_counter_RNO_0_3_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__27996),
            .in2(N__27949),
            .in3(N__26461),
            .lcout(\ws2812.rgb_counter_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\ws2812.un1_rgb_counter_cry_2 ),
            .carryout(\ws2812.un1_rgb_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_0_3_LC_12_8_4 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_3_LC_12_8_4 .SEQ_MODE=4'b1011;
    defparam \ws2812.rgb_counter_0_3_LC_12_8_4 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \ws2812.rgb_counter_0_3_LC_12_8_4  (
            .in0(N__27711),
            .in1(N__27861),
            .in2(N__26755),
            .in3(N__26692),
            .lcout(\ws2812.rgb_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27509),
            .ce(),
            .sr(N__27132));
    defparam \ws2812.rgb_counter_0_RNIP62Q_3_LC_12_9_0 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_RNIP62Q_3_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_0_RNIP62Q_3_LC_12_9_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ws2812.rgb_counter_0_RNIP62Q_3_LC_12_9_0  (
            .in0(N__26689),
            .in1(N__26745),
            .in2(N__26617),
            .in3(N__28108),
            .lcout(),
            .ltout(\ws2812.rgb_data_pmux_10_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIOLAI1_2_LC_12_9_1 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIOLAI1_2_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIOLAI1_2_LC_12_9_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ws2812.rgb_counter_RNIOLAI1_2_LC_12_9_1  (
            .in0(N__28109),
            .in1(N__26683),
            .in2(N__26677),
            .in3(N__26674),
            .lcout(\ws2812.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_0_RNIR82Q_3_LC_12_9_6 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_RNIR82Q_3_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_0_RNIR82Q_3_LC_12_9_6 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \ws2812.rgb_counter_0_RNIR82Q_3_LC_12_9_6  (
            .in0(N__26632),
            .in1(N__26659),
            .in2(N__28122),
            .in3(N__26744),
            .lcout(\ws2812.rgb_data_pmux_6_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_out_2_LC_12_9_7 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_2_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_2_LC_12_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_2_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26647),
            .lcout(rgb_data_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27515),
            .ce(N__27195),
            .sr(N__27136));
    defparam \sb_translator_1.rgb_data_out_17_LC_12_10_1 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_17_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_17_LC_12_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sb_translator_1.rgb_data_out_17_LC_12_10_1  (
            .in0(N__26626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_data_out_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27517),
            .ce(N__27192),
            .sr(N__27138));
    defparam \sb_translator_1.rgb_data_out_23_LC_12_10_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_23_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_23_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_23_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26608),
            .lcout(rgb_data_out_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27517),
            .ce(N__27192),
            .sr(N__27138));
    defparam \sb_translator_1.rgb_data_out_14_LC_12_10_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_14_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_14_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_14_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26599),
            .lcout(rgb_data_out_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27517),
            .ce(N__27192),
            .sr(N__27138));
    defparam \sb_translator_1.rgb_data_out_22_LC_12_10_7 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_22_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_22_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_22_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26914),
            .lcout(rgb_data_out_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27517),
            .ce(N__27192),
            .sr(N__27138));
    defparam \ws2812.state_0_LC_13_6_0 .C_ON=1'b0;
    defparam \ws2812.state_0_LC_13_6_0 .SEQ_MODE=4'b1011;
    defparam \ws2812.state_0_LC_13_6_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ws2812.state_0_LC_13_6_0  (
            .in0(N__27562),
            .in1(N__27679),
            .in2(_gnd_net_),
            .in3(N__26904),
            .lcout(\ws2812.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27506),
            .ce(),
            .sr(N__27129));
    defparam \ws2812.rgb_counter_0_RNITA2Q_3_LC_13_7_0 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_0_RNITA2Q_3_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_0_RNITA2Q_3_LC_13_7_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ws2812.rgb_counter_0_RNITA2Q_3_LC_13_7_0  (
            .in0(N__26800),
            .in1(N__26749),
            .in2(N__26782),
            .in3(N__28112),
            .lcout(),
            .ltout(\ws2812.rgb_data_pmux_13_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI0UAI1_2_LC_13_7_1 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI0UAI1_2_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI0UAI1_2_LC_13_7_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ws2812.rgb_counter_RNI0UAI1_2_LC_13_7_1  (
            .in0(N__28113),
            .in1(N__26830),
            .in2(N__26821),
            .in3(N__26761),
            .lcout(\ws2812.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_out_3_LC_13_7_2 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_3_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_3_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_3_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26812),
            .lcout(rgb_data_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27510),
            .ce(N__27197),
            .sr(N__27133));
    defparam \sb_translator_1.rgb_data_out_19_LC_13_7_3 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_19_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_19_LC_13_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_19_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26794),
            .lcout(rgb_data_out_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27510),
            .ce(N__27197),
            .sr(N__27133));
    defparam \sb_translator_1.rgb_data_out_7_LC_13_7_4 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_7_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_7_LC_13_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_7_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26773),
            .lcout(rgb_data_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27510),
            .ce(N__27197),
            .sr(N__27133));
    defparam \ws2812.rgb_counter_RNIRMNJ1_3_LC_13_7_7 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIRMNJ1_3_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIRMNJ1_3_LC_13_7_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ws2812.rgb_counter_RNIRMNJ1_3_LC_13_7_7  (
            .in0(N__26750),
            .in1(N__27995),
            .in2(N__28132),
            .in3(N__28034),
            .lcout(\ws2812.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNISPAI1_2_LC_13_8_0 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNISPAI1_2_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNISPAI1_2_LC_13_8_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ws2812.rgb_counter_RNISPAI1_2_LC_13_8_0  (
            .in0(N__27526),
            .in1(N__28110),
            .in2(N__26719),
            .in3(N__26707),
            .lcout(\ws2812.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNIGEUO_0_LC_13_8_2 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNIGEUO_0_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNIGEUO_0_LC_13_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ws2812.rgb_counter_RNIGEUO_0_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__27935),
            .in2(_gnd_net_),
            .in3(N__28111),
            .lcout(\ws2812.rgb_counter_0_sqmuxa_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI2AOD3_2_LC_13_8_3 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI2AOD3_2_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI2AOD3_2_LC_13_8_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \ws2812.rgb_counter_RNI2AOD3_2_LC_13_8_3  (
            .in0(N__27858),
            .in1(_gnd_net_),
            .in2(N__27742),
            .in3(N__28123),
            .lcout(\ws2812.rgb_counter_RNI2AOD3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI19OD3_1_LC_13_8_4 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI19OD3_1_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI19OD3_1_LC_13_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ws2812.rgb_counter_RNI19OD3_1_LC_13_8_4  (
            .in0(N__28039),
            .in1(N__27701),
            .in2(_gnd_net_),
            .in3(N__27857),
            .lcout(\ws2812.rgb_counter_RNI19OD3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.rgb_counter_RNI3BOD3_3_LC_13_8_5 .C_ON=1'b0;
    defparam \ws2812.rgb_counter_RNI3BOD3_3_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \ws2812.rgb_counter_RNI3BOD3_3_LC_13_8_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \ws2812.rgb_counter_RNI3BOD3_3_LC_13_8_5  (
            .in0(N__27859),
            .in1(N__27997),
            .in2(N__27743),
            .in3(_gnd_net_),
            .lcout(\ws2812.rgb_counter_RNI3BOD3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.un1_rgb_counter_cry_0_c_RNO_LC_13_8_6 .C_ON=1'b0;
    defparam \ws2812.un1_rgb_counter_cry_0_c_RNO_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \ws2812.un1_rgb_counter_cry_0_c_RNO_LC_13_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ws2812.un1_rgb_counter_cry_0_c_RNO_LC_13_8_6  (
            .in0(N__27940),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__27700),
            .lcout(\ws2812.un1_rgb_counter_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ws2812.state_RNIELS35_0_LC_13_8_7 .C_ON=1'b0;
    defparam \ws2812.state_RNIELS35_0_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \ws2812.state_RNIELS35_0_LC_13_8_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \ws2812.state_RNIELS35_0_LC_13_8_7  (
            .in0(N__27860),
            .in1(N__27787),
            .in2(N__27744),
            .in3(N__27588),
            .lcout(\ws2812.state_RNIELS35Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sb_translator_1.rgb_data_out_6_LC_13_9_5 .C_ON=1'b0;
    defparam \sb_translator_1.rgb_data_out_6_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \sb_translator_1.rgb_data_out_6_LC_13_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sb_translator_1.rgb_data_out_6_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27535),
            .lcout(rgb_data_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__27518),
            .ce(N__27196),
            .sr(N__27139));
endmodule // top
